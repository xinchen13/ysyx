//Generate the verilog at 2024-08-23T20:33:26
module alu1 (
clk,
a,
b,
ctrl,
result
);

input clk ;
input [31:0] a ;
input [31:0] b ;
input [3:0] ctrl ;
output [31:0] result ;

wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire _133_ ;
wire _134_ ;
wire _135_ ;
wire _136_ ;
wire _137_ ;
wire _138_ ;
wire _139_ ;
wire _140_ ;
wire _141_ ;
wire _142_ ;
wire _143_ ;
wire _144_ ;
wire _145_ ;
wire _146_ ;
wire _147_ ;
wire _148_ ;
wire _149_ ;
wire _150_ ;
wire _151_ ;
wire _152_ ;
wire _153_ ;
wire _154_ ;
wire _155_ ;
wire _156_ ;
wire _157_ ;
wire _158_ ;
wire _159_ ;
wire _160_ ;
wire _161_ ;
wire _162_ ;
wire _163_ ;
wire _164_ ;
wire _165_ ;
wire _166_ ;
wire _167_ ;
wire _168_ ;
wire _169_ ;
wire _170_ ;
wire _171_ ;
wire _172_ ;
wire _173_ ;
wire _174_ ;
wire _175_ ;
wire _176_ ;
wire _177_ ;
wire _178_ ;
wire _179_ ;
wire _180_ ;
wire _181_ ;
wire _182_ ;
wire _183_ ;
wire _184_ ;
wire _185_ ;
wire _186_ ;
wire _187_ ;
wire _188_ ;
wire _189_ ;
wire _190_ ;
wire _191_ ;
wire _192_ ;
wire _193_ ;
wire _194_ ;
wire _195_ ;
wire _196_ ;
wire _197_ ;
wire _198_ ;
wire _199_ ;
wire _200_ ;
wire _201_ ;
wire _202_ ;
wire _203_ ;
wire _204_ ;
wire _205_ ;
wire _206_ ;
wire _207_ ;
wire _208_ ;
wire _209_ ;
wire _210_ ;
wire _211_ ;
wire _212_ ;
wire _213_ ;
wire _214_ ;
wire _215_ ;
wire _216_ ;
wire _217_ ;
wire _218_ ;
wire _219_ ;
wire _220_ ;
wire _221_ ;
wire _222_ ;
wire _223_ ;
wire _224_ ;
wire _225_ ;
wire _226_ ;
wire _227_ ;
wire _228_ ;
wire _229_ ;
wire _230_ ;
wire _231_ ;
wire _232_ ;
wire _233_ ;
wire _234_ ;
wire _235_ ;
wire _236_ ;
wire _237_ ;
wire _238_ ;
wire _239_ ;
wire _240_ ;
wire _241_ ;
wire _242_ ;
wire _243_ ;
wire _244_ ;
wire _245_ ;
wire _246_ ;
wire _247_ ;
wire _248_ ;
wire _249_ ;
wire _250_ ;
wire _251_ ;
wire _252_ ;
wire _253_ ;
wire _254_ ;
wire _255_ ;
wire _256_ ;
wire _257_ ;
wire _258_ ;
wire _259_ ;
wire _260_ ;
wire _261_ ;
wire _262_ ;
wire _263_ ;
wire _264_ ;
wire _265_ ;
wire _266_ ;
wire _267_ ;
wire _268_ ;
wire _269_ ;
wire _270_ ;
wire _271_ ;
wire _272_ ;
wire _273_ ;
wire _274_ ;
wire _275_ ;
wire _276_ ;
wire _277_ ;
wire _278_ ;
wire _279_ ;
wire _280_ ;
wire _281_ ;
wire _282_ ;
wire _283_ ;
wire _284_ ;
wire _285_ ;
wire _286_ ;
wire _287_ ;
wire _288_ ;
wire _289_ ;
wire _290_ ;
wire _291_ ;
wire _292_ ;
wire _293_ ;
wire _294_ ;
wire _295_ ;
wire _296_ ;
wire _297_ ;
wire _298_ ;
wire _299_ ;
wire _300_ ;
wire _301_ ;
wire _302_ ;
wire _303_ ;
wire _304_ ;
wire _305_ ;
wire _306_ ;
wire _307_ ;
wire _308_ ;
wire _309_ ;
wire _310_ ;
wire _311_ ;
wire _312_ ;
wire _313_ ;
wire _314_ ;
wire _315_ ;
wire _316_ ;
wire _317_ ;
wire _318_ ;
wire _319_ ;
wire _320_ ;
wire _321_ ;
wire _322_ ;
wire _323_ ;
wire _324_ ;
wire _325_ ;
wire _326_ ;
wire _327_ ;
wire _328_ ;
wire _329_ ;
wire _330_ ;
wire _331_ ;
wire _332_ ;
wire _333_ ;
wire _334_ ;
wire _335_ ;
wire _336_ ;
wire _337_ ;
wire _338_ ;
wire _339_ ;
wire _340_ ;
wire _341_ ;
wire _342_ ;
wire _343_ ;
wire _344_ ;
wire _345_ ;
wire _346_ ;
wire _347_ ;
wire _348_ ;
wire _349_ ;
wire _350_ ;
wire _351_ ;
wire _352_ ;
wire _353_ ;
wire _354_ ;
wire _355_ ;
wire _356_ ;
wire _357_ ;
wire _358_ ;
wire _359_ ;
wire _360_ ;
wire _361_ ;
wire _362_ ;
wire _363_ ;
wire _364_ ;
wire _365_ ;
wire _366_ ;
wire _367_ ;
wire _368_ ;
wire _369_ ;
wire _370_ ;
wire _371_ ;
wire _372_ ;
wire _373_ ;
wire _374_ ;
wire _375_ ;
wire _376_ ;
wire _377_ ;
wire _378_ ;
wire _379_ ;
wire _380_ ;
wire _381_ ;
wire _382_ ;
wire _383_ ;
wire _384_ ;
wire _385_ ;
wire _386_ ;
wire _387_ ;
wire _388_ ;
wire _389_ ;
wire _390_ ;
wire _391_ ;
wire _392_ ;
wire _393_ ;
wire _394_ ;
wire _395_ ;
wire _396_ ;
wire _397_ ;
wire _398_ ;
wire _399_ ;
wire _400_ ;
wire _401_ ;
wire _402_ ;
wire _403_ ;
wire _404_ ;
wire _405_ ;
wire _406_ ;
wire _407_ ;
wire _408_ ;
wire _409_ ;
wire _410_ ;
wire _411_ ;
wire _412_ ;
wire _413_ ;
wire _414_ ;
wire _415_ ;
wire _416_ ;
wire _417_ ;
wire _418_ ;
wire _419_ ;
wire _420_ ;
wire _421_ ;
wire _422_ ;
wire _423_ ;
wire _424_ ;
wire _425_ ;
wire _426_ ;
wire _427_ ;
wire _428_ ;
wire _429_ ;
wire _430_ ;
wire _431_ ;
wire _432_ ;
wire _433_ ;
wire _434_ ;
wire _435_ ;
wire _436_ ;
wire _437_ ;
wire _438_ ;
wire _439_ ;
wire _440_ ;
wire _441_ ;
wire [31:0] b ;
wire [31:0] a ;
wire [3:0] ctrl ;
wire [31:0] result ;


XNOR2_X2 _442_ ( .A(_005_ ), .B(_037_ ), .ZN(_068_ ) );
XNOR2_X2 _443_ ( .A(_006_ ), .B(_038_ ), .ZN(_069_ ) );
AND2_X4 _444_ ( .A1(_068_ ), .A2(_069_ ), .ZN(_070_ ) );
XNOR2_X2 _445_ ( .A(_004_ ), .B(_036_ ), .ZN(_071_ ) );
XNOR2_X2 _446_ ( .A(_003_ ), .B(_035_ ), .ZN(_072_ ) );
AND2_X2 _447_ ( .A1(_071_ ), .A2(_072_ ), .ZN(_073_ ) );
AND2_X4 _448_ ( .A1(_070_ ), .A2(_073_ ), .ZN(_074_ ) );
XNOR2_X2 _449_ ( .A(_001_ ), .B(_033_ ), .ZN(_075_ ) );
XNOR2_X2 _450_ ( .A(_002_ ), .B(_034_ ), .ZN(_076_ ) );
AND2_X1 _451_ ( .A1(_075_ ), .A2(_076_ ), .ZN(_077_ ) );
XNOR2_X2 _452_ ( .A(_031_ ), .B(_063_ ), .ZN(_078_ ) );
XNOR2_X1 _453_ ( .A(_030_ ), .B(_062_ ), .ZN(_079_ ) );
AND3_X2 _454_ ( .A1(_077_ ), .A2(_078_ ), .A3(_079_ ), .ZN(_080_ ) );
XNOR2_X2 _455_ ( .A(_028_ ), .B(_060_ ), .ZN(_081_ ) );
XNOR2_X2 _456_ ( .A(_029_ ), .B(_061_ ), .ZN(_082_ ) );
AND2_X1 _457_ ( .A1(_081_ ), .A2(_082_ ), .ZN(_083_ ) );
XNOR2_X1 _458_ ( .A(_026_ ), .B(_058_ ), .ZN(_084_ ) );
XNOR2_X2 _459_ ( .A(_027_ ), .B(_059_ ), .ZN(_085_ ) );
AND3_X1 _460_ ( .A1(_083_ ), .A2(_084_ ), .A3(_085_ ), .ZN(_086_ ) );
XNOR2_X2 _461_ ( .A(_022_ ), .B(_054_ ), .ZN(_087_ ) );
XNOR2_X2 _462_ ( .A(_025_ ), .B(_057_ ), .ZN(_088_ ) );
XNOR2_X2 _463_ ( .A(_011_ ), .B(_043_ ), .ZN(_089_ ) );
XNOR2_X1 _464_ ( .A(_032_ ), .B(_000_ ), .ZN(_090_ ) );
AND4_X1 _465_ ( .A1(_087_ ), .A2(_088_ ), .A3(_089_ ), .A4(_090_ ), .ZN(_091_ ) );
AND4_X1 _466_ ( .A1(_074_ ), .A2(_080_ ), .A3(_086_ ), .A4(_091_ ), .ZN(_092_ ) );
XNOR2_X1 _467_ ( .A(_009_ ), .B(_041_ ), .ZN(_093_ ) );
XNOR2_X1 _468_ ( .A(_010_ ), .B(_042_ ), .ZN(_094_ ) );
AND2_X1 _469_ ( .A1(_093_ ), .A2(_094_ ), .ZN(_095_ ) );
XNOR2_X1 _470_ ( .A(_008_ ), .B(_040_ ), .ZN(_096_ ) );
XNOR2_X1 _471_ ( .A(_007_ ), .B(_039_ ), .ZN(_097_ ) );
AND3_X1 _472_ ( .A1(_095_ ), .A2(_096_ ), .A3(_097_ ), .ZN(_098_ ) );
XNOR2_X1 _473_ ( .A(_012_ ), .B(_044_ ), .ZN(_099_ ) );
XNOR2_X1 _474_ ( .A(_013_ ), .B(_045_ ), .ZN(_100_ ) );
AND2_X1 _475_ ( .A1(_099_ ), .A2(_100_ ), .ZN(_101_ ) );
XNOR2_X1 _476_ ( .A(_014_ ), .B(_046_ ), .ZN(_102_ ) );
XNOR2_X1 _477_ ( .A(_015_ ), .B(_047_ ), .ZN(_103_ ) );
AND2_X1 _478_ ( .A1(_102_ ), .A2(_103_ ), .ZN(_104_ ) );
AND2_X1 _479_ ( .A1(_101_ ), .A2(_104_ ), .ZN(_105_ ) );
AND2_X1 _480_ ( .A1(_098_ ), .A2(_105_ ), .ZN(_106_ ) );
XNOR2_X1 _481_ ( .A(_023_ ), .B(_055_ ), .ZN(_107_ ) );
XNOR2_X1 _482_ ( .A(_024_ ), .B(_056_ ), .ZN(_108_ ) );
AND2_X1 _483_ ( .A1(_107_ ), .A2(_108_ ), .ZN(_109_ ) );
XNOR2_X1 _484_ ( .A(_020_ ), .B(_052_ ), .ZN(_110_ ) );
XNOR2_X1 _485_ ( .A(_021_ ), .B(_053_ ), .ZN(_111_ ) );
AND3_X1 _486_ ( .A1(_109_ ), .A2(_110_ ), .A3(_111_ ), .ZN(_112_ ) );
XNOR2_X1 _487_ ( .A(_018_ ), .B(_050_ ), .ZN(_113_ ) );
XNOR2_X1 _488_ ( .A(_019_ ), .B(_051_ ), .ZN(_114_ ) );
AND2_X1 _489_ ( .A1(_113_ ), .A2(_114_ ), .ZN(_115_ ) );
XNOR2_X1 _490_ ( .A(_017_ ), .B(_049_ ), .ZN(_116_ ) );
XNOR2_X1 _491_ ( .A(_016_ ), .B(_048_ ), .ZN(_117_ ) );
AND3_X1 _492_ ( .A1(_115_ ), .A2(_116_ ), .A3(_117_ ), .ZN(_118_ ) );
AND2_X1 _493_ ( .A1(_112_ ), .A2(_118_ ), .ZN(_119_ ) );
NAND3_X1 _494_ ( .A1(_092_ ), .A2(_106_ ), .A3(_119_ ), .ZN(_120_ ) );
NOR2_X1 _495_ ( .A1(_064_ ), .A2(_066_ ), .ZN(_121_ ) );
NAND3_X1 _496_ ( .A1(_120_ ), .A2(_067_ ), .A3(_121_ ), .ZN(_122_ ) );
INV_X1 _497_ ( .A(_020_ ), .ZN(_123_ ) );
AND3_X1 _498_ ( .A1(_111_ ), .A2(_123_ ), .A3(_052_ ), .ZN(_124_ ) );
INV_X1 _499_ ( .A(_053_ ), .ZN(_125_ ) );
NOR2_X1 _500_ ( .A1(_125_ ), .A2(_021_ ), .ZN(_126_ ) );
OAI21_X1 _501_ ( .A(_109_ ), .B1(_124_ ), .B2(_126_ ), .ZN(_127_ ) );
INV_X1 _502_ ( .A(_047_ ), .ZN(_128_ ) );
NOR2_X1 _503_ ( .A1(_128_ ), .A2(_015_ ), .ZN(_129_ ) );
INV_X1 _504_ ( .A(_129_ ), .ZN(_130_ ) );
INV_X1 _505_ ( .A(_045_ ), .ZN(_131_ ) );
AND2_X1 _506_ ( .A1(_131_ ), .A2(_013_ ), .ZN(_132_ ) );
NOR2_X1 _507_ ( .A1(_131_ ), .A2(_013_ ), .ZN(_133_ ) );
INV_X1 _508_ ( .A(_044_ ), .ZN(_134_ ) );
NOR4_X1 _509_ ( .A1(_132_ ), .A2(_133_ ), .A3(_012_ ), .A4(_134_ ), .ZN(_135_ ) );
OAI21_X1 _510_ ( .A(_104_ ), .B1(_135_ ), .B2(_133_ ), .ZN(_136_ ) );
INV_X1 _511_ ( .A(_008_ ), .ZN(_137_ ) );
AND2_X1 _512_ ( .A1(_137_ ), .A2(_040_ ), .ZN(_138_ ) );
NOR2_X1 _513_ ( .A1(_137_ ), .A2(_040_ ), .ZN(_139_ ) );
INV_X1 _514_ ( .A(_039_ ), .ZN(_140_ ) );
NOR4_X1 _515_ ( .A1(_138_ ), .A2(_139_ ), .A3(_007_ ), .A4(_140_ ), .ZN(_141_ ) );
OAI21_X1 _516_ ( .A(_095_ ), .B1(_141_ ), .B2(_138_ ), .ZN(_142_ ) );
INV_X1 _517_ ( .A(_042_ ), .ZN(_143_ ) );
NOR2_X1 _518_ ( .A1(_143_ ), .A2(_010_ ), .ZN(_144_ ) );
INV_X1 _519_ ( .A(_144_ ), .ZN(_145_ ) );
INV_X1 _520_ ( .A(_009_ ), .ZN(_146_ ) );
NAND3_X1 _521_ ( .A1(_094_ ), .A2(_146_ ), .A3(_041_ ), .ZN(_147_ ) );
AND3_X1 _522_ ( .A1(_142_ ), .A2(_145_ ), .A3(_147_ ), .ZN(_148_ ) );
INV_X1 _523_ ( .A(_105_ ), .ZN(_149_ ) );
OAI211_X2 _524_ ( .A(_130_ ), .B(_136_ ), .C1(_148_ ), .C2(_149_ ), .ZN(_150_ ) );
INV_X1 _525_ ( .A(_046_ ), .ZN(_151_ ) );
AOI211_X4 _526_ ( .A(_014_ ), .B(_151_ ), .C1(_015_ ), .C2(_128_ ), .ZN(_152_ ) );
OAI21_X1 _527_ ( .A(_119_ ), .B1(_150_ ), .B2(_152_ ), .ZN(_153_ ) );
INV_X1 _528_ ( .A(_023_ ), .ZN(_154_ ) );
AND2_X1 _529_ ( .A1(_154_ ), .A2(_055_ ), .ZN(_155_ ) );
INV_X1 _530_ ( .A(_024_ ), .ZN(_156_ ) );
OAI21_X1 _531_ ( .A(_155_ ), .B1(_156_ ), .B2(_056_ ), .ZN(_157_ ) );
INV_X1 _532_ ( .A(_115_ ), .ZN(_158_ ) );
INV_X1 _533_ ( .A(_017_ ), .ZN(_159_ ) );
AND2_X1 _534_ ( .A1(_159_ ), .A2(_049_ ), .ZN(_160_ ) );
INV_X1 _535_ ( .A(_160_ ), .ZN(_161_ ) );
INV_X1 _536_ ( .A(_048_ ), .ZN(_162_ ) );
NOR2_X1 _537_ ( .A1(_162_ ), .A2(_016_ ), .ZN(_163_ ) );
NAND2_X1 _538_ ( .A1(_116_ ), .A2(_163_ ), .ZN(_164_ ) );
AOI21_X1 _539_ ( .A(_158_ ), .B1(_161_ ), .B2(_164_ ), .ZN(_165_ ) );
INV_X1 _540_ ( .A(_019_ ), .ZN(_166_ ) );
AND2_X1 _541_ ( .A1(_166_ ), .A2(_051_ ), .ZN(_167_ ) );
INV_X1 _542_ ( .A(_018_ ), .ZN(_168_ ) );
AND3_X1 _543_ ( .A1(_114_ ), .A2(_168_ ), .A3(_050_ ), .ZN(_169_ ) );
OR3_X1 _544_ ( .A1(_165_ ), .A2(_167_ ), .A3(_169_ ), .ZN(_170_ ) );
AOI22_X1 _545_ ( .A1(_170_ ), .A2(_112_ ), .B1(_156_ ), .B2(_056_ ), .ZN(_171_ ) );
AND4_X1 _546_ ( .A1(_127_ ), .A2(_153_ ), .A3(_157_ ), .A4(_171_ ), .ZN(_172_ ) );
AND2_X1 _547_ ( .A1(_119_ ), .A2(_106_ ), .ZN(_173_ ) );
INV_X4 _548_ ( .A(_062_ ), .ZN(_174_ ) );
NOR2_X1 _549_ ( .A1(_174_ ), .A2(_030_ ), .ZN(_175_ ) );
AND2_X1 _550_ ( .A1(_078_ ), .A2(_175_ ), .ZN(_176_ ) );
INV_X2 _551_ ( .A(_031_ ), .ZN(_177_ ) );
AND2_X1 _552_ ( .A1(_177_ ), .A2(_063_ ), .ZN(_178_ ) );
OAI21_X1 _553_ ( .A(_077_ ), .B1(_176_ ), .B2(_178_ ), .ZN(_179_ ) );
INV_X2 _554_ ( .A(_001_ ), .ZN(_180_ ) );
INV_X1 _555_ ( .A(_002_ ), .ZN(_181_ ) );
OAI211_X2 _556_ ( .A(_180_ ), .B(_033_ ), .C1(_181_ ), .C2(_034_ ), .ZN(_182_ ) );
NAND2_X1 _557_ ( .A1(_179_ ), .A2(_182_ ), .ZN(_183_ ) );
AOI21_X1 _558_ ( .A(_183_ ), .B1(_181_ ), .B2(_034_ ), .ZN(_184_ ) );
INV_X2 _559_ ( .A(_074_ ), .ZN(_185_ ) );
OR2_X1 _560_ ( .A1(_184_ ), .A2(_185_ ), .ZN(_186_ ) );
INV_X1 _561_ ( .A(_006_ ), .ZN(_187_ ) );
AND2_X1 _562_ ( .A1(_187_ ), .A2(_038_ ), .ZN(_188_ ) );
INV_X1 _563_ ( .A(_188_ ), .ZN(_189_ ) );
INV_X16 _564_ ( .A(_035_ ), .ZN(_190_ ) );
NOR2_X1 _565_ ( .A1(_190_ ), .A2(_003_ ), .ZN(_191_ ) );
AND2_X1 _566_ ( .A1(_071_ ), .A2(_191_ ), .ZN(_192_ ) );
INV_X1 _567_ ( .A(_004_ ), .ZN(_193_ ) );
AND2_X1 _568_ ( .A1(_193_ ), .A2(_036_ ), .ZN(_194_ ) );
OAI21_X1 _569_ ( .A(_070_ ), .B1(_192_ ), .B2(_194_ ), .ZN(_195_ ) );
NOR2_X1 _570_ ( .A1(_187_ ), .A2(_038_ ), .ZN(_196_ ) );
INV_X1 _571_ ( .A(_037_ ), .ZN(_197_ ) );
OR4_X1 _572_ ( .A1(_005_ ), .A2(_188_ ), .A3(_196_ ), .A4(_197_ ), .ZN(_198_ ) );
NAND4_X1 _573_ ( .A1(_186_ ), .A2(_189_ ), .A3(_195_ ), .A4(_198_ ), .ZN(_199_ ) );
AND2_X1 _574_ ( .A1(_080_ ), .A2(_074_ ), .ZN(_200_ ) );
INV_X1 _575_ ( .A(_200_ ), .ZN(_201_ ) );
INV_X16 _576_ ( .A(_000_ ), .ZN(_202_ ) );
INV_X1 _577_ ( .A(_011_ ), .ZN(_203_ ) );
AOI211_X4 _578_ ( .A(_032_ ), .B(_202_ ), .C1(_203_ ), .C2(_043_ ), .ZN(_204_ ) );
INV_X1 _579_ ( .A(_087_ ), .ZN(_205_ ) );
INV_X1 _580_ ( .A(_088_ ), .ZN(_206_ ) );
NOR2_X1 _581_ ( .A1(_203_ ), .A2(_043_ ), .ZN(_207_ ) );
NOR4_X1 _582_ ( .A1(_204_ ), .A2(_205_ ), .A3(_206_ ), .A4(_207_ ), .ZN(_208_ ) );
INV_X1 _583_ ( .A(_022_ ), .ZN(_209_ ) );
NAND3_X1 _584_ ( .A1(_088_ ), .A2(_209_ ), .A3(_054_ ), .ZN(_210_ ) );
INV_X1 _585_ ( .A(_057_ ), .ZN(_211_ ) );
NOR2_X1 _586_ ( .A1(_211_ ), .A2(_025_ ), .ZN(_212_ ) );
INV_X1 _587_ ( .A(_212_ ), .ZN(_213_ ) );
NAND2_X1 _588_ ( .A1(_210_ ), .A2(_213_ ), .ZN(_214_ ) );
OAI21_X1 _589_ ( .A(_086_ ), .B1(_208_ ), .B2(_214_ ), .ZN(_215_ ) );
INV_X1 _590_ ( .A(_058_ ), .ZN(_216_ ) );
NOR2_X1 _591_ ( .A1(_216_ ), .A2(_026_ ), .ZN(_217_ ) );
AND2_X1 _592_ ( .A1(_085_ ), .A2(_217_ ), .ZN(_218_ ) );
INV_X2 _593_ ( .A(_059_ ), .ZN(_219_ ) );
NOR2_X1 _594_ ( .A1(_219_ ), .A2(_027_ ), .ZN(_220_ ) );
OAI21_X1 _595_ ( .A(_083_ ), .B1(_218_ ), .B2(_220_ ), .ZN(_221_ ) );
INV_X1 _596_ ( .A(_061_ ), .ZN(_222_ ) );
NOR2_X1 _597_ ( .A1(_222_ ), .A2(_029_ ), .ZN(_223_ ) );
INV_X1 _598_ ( .A(_028_ ), .ZN(_224_ ) );
AND2_X1 _599_ ( .A1(_224_ ), .A2(_060_ ), .ZN(_225_ ) );
AOI21_X1 _600_ ( .A(_223_ ), .B1(_082_ ), .B2(_225_ ), .ZN(_226_ ) );
AND2_X1 _601_ ( .A1(_221_ ), .A2(_226_ ), .ZN(_227_ ) );
AOI21_X1 _602_ ( .A(_201_ ), .B1(_215_ ), .B2(_227_ ), .ZN(_228_ ) );
OAI21_X1 _603_ ( .A(_173_ ), .B1(_199_ ), .B2(_228_ ), .ZN(_229_ ) );
AOI21_X1 _604_ ( .A(_122_ ), .B1(_172_ ), .B2(_229_ ), .ZN(_230_ ) );
NAND2_X1 _605_ ( .A1(_230_ ), .A2(_065_ ), .ZN(_231_ ) );
INV_X1 _606_ ( .A(_121_ ), .ZN(_232_ ) );
NOR2_X1 _607_ ( .A1(_232_ ), .A2(_065_ ), .ZN(_233_ ) );
INV_X1 _608_ ( .A(_233_ ), .ZN(_234_ ) );
BUF_X4 _609_ ( .A(_234_ ), .Z(_235_ ) );
OAI21_X1 _610_ ( .A(_231_ ), .B1(_090_ ), .B2(_235_ ), .ZN(_410_ ) );
AND2_X1 _611_ ( .A1(_202_ ), .A2(_032_ ), .ZN(_236_ ) );
INV_X1 _612_ ( .A(_236_ ), .ZN(_237_ ) );
OAI21_X1 _613_ ( .A(_233_ ), .B1(_237_ ), .B2(_089_ ), .ZN(_238_ ) );
AOI21_X1 _614_ ( .A(_238_ ), .B1(_089_ ), .B2(_237_ ), .ZN(_421_ ) );
NAND2_X1 _615_ ( .A1(_237_ ), .A2(_089_ ), .ZN(_239_ ) );
INV_X1 _616_ ( .A(_207_ ), .ZN(_240_ ) );
AND3_X1 _617_ ( .A1(_239_ ), .A2(_205_ ), .A3(_240_ ), .ZN(_241_ ) );
AOI21_X1 _618_ ( .A(_205_ ), .B1(_239_ ), .B2(_240_ ), .ZN(_242_ ) );
NOR3_X1 _619_ ( .A1(_241_ ), .A2(_242_ ), .A3(_234_ ), .ZN(_432_ ) );
NOR2_X2 _620_ ( .A1(_209_ ), .A2(_054_ ), .ZN(_243_ ) );
OR3_X1 _621_ ( .A1(_242_ ), .A2(_243_ ), .A3(_088_ ), .ZN(_244_ ) );
CLKBUF_X2 _622_ ( .A(_233_ ), .Z(_245_ ) );
OAI21_X1 _623_ ( .A(_088_ ), .B1(_242_ ), .B2(_243_ ), .ZN(_246_ ) );
AND3_X1 _624_ ( .A1(_244_ ), .A2(_245_ ), .A3(_246_ ), .ZN(_435_ ) );
AND2_X2 _625_ ( .A1(_088_ ), .A2(_243_ ), .ZN(_247_ ) );
AOI21_X2 _626_ ( .A(_247_ ), .B1(_025_ ), .B2(_211_ ), .ZN(_248_ ) );
INV_X1 _627_ ( .A(_248_ ), .ZN(_249_ ) );
AOI211_X2 _628_ ( .A(_205_ ), .B(_206_ ), .C1(_239_ ), .C2(_240_ ), .ZN(_250_ ) );
NOR2_X2 _629_ ( .A1(_249_ ), .A2(_250_ ), .ZN(_251_ ) );
INV_X2 _630_ ( .A(_251_ ), .ZN(_252_ ) );
OAI21_X1 _631_ ( .A(_245_ ), .B1(_252_ ), .B2(_084_ ), .ZN(_253_ ) );
INV_X1 _632_ ( .A(_084_ ), .ZN(_254_ ) );
NOR2_X1 _633_ ( .A1(_251_ ), .A2(_254_ ), .ZN(_255_ ) );
NOR2_X1 _634_ ( .A1(_253_ ), .A2(_255_ ), .ZN(_436_ ) );
AND2_X1 _635_ ( .A1(_216_ ), .A2(_026_ ), .ZN(_256_ ) );
OR3_X1 _636_ ( .A1(_255_ ), .A2(_256_ ), .A3(_085_ ), .ZN(_257_ ) );
OAI21_X1 _637_ ( .A(_085_ ), .B1(_255_ ), .B2(_256_ ), .ZN(_258_ ) );
AND3_X1 _638_ ( .A1(_257_ ), .A2(_245_ ), .A3(_258_ ), .ZN(_437_ ) );
AND2_X4 _639_ ( .A1(_219_ ), .A2(_027_ ), .ZN(_259_ ) );
NOR4_X1 _640_ ( .A1(_251_ ), .A2(_220_ ), .A3(_259_ ), .A4(_254_ ), .ZN(_260_ ) );
AOI21_X1 _641_ ( .A(_259_ ), .B1(_085_ ), .B2(_256_ ), .ZN(_261_ ) );
INV_X1 _642_ ( .A(_261_ ), .ZN(_262_ ) );
NOR2_X1 _643_ ( .A1(_260_ ), .A2(_262_ ), .ZN(_263_ ) );
INV_X1 _644_ ( .A(_081_ ), .ZN(_264_ ) );
NOR2_X1 _645_ ( .A1(_263_ ), .A2(_264_ ), .ZN(_265_ ) );
NOR3_X1 _646_ ( .A1(_260_ ), .A2(_081_ ), .A3(_262_ ), .ZN(_266_ ) );
NOR3_X1 _647_ ( .A1(_265_ ), .A2(_235_ ), .A3(_266_ ), .ZN(_438_ ) );
NOR2_X1 _648_ ( .A1(_224_ ), .A2(_060_ ), .ZN(_267_ ) );
OR3_X1 _649_ ( .A1(_265_ ), .A2(_267_ ), .A3(_082_ ), .ZN(_268_ ) );
OAI21_X1 _650_ ( .A(_082_ ), .B1(_265_ ), .B2(_267_ ), .ZN(_269_ ) );
AND3_X1 _651_ ( .A1(_268_ ), .A2(_245_ ), .A3(_269_ ), .ZN(_439_ ) );
AND2_X4 _652_ ( .A1(_252_ ), .A2(_086_ ), .ZN(_270_ ) );
AND2_X2 _653_ ( .A1(_082_ ), .A2(_267_ ), .ZN(_271_ ) );
AOI221_X1 _654_ ( .A(_271_ ), .B1(_029_ ), .B2(_222_ ), .C1(_262_ ), .C2(_083_ ), .ZN(_272_ ) );
INV_X2 _655_ ( .A(_272_ ), .ZN(_273_ ) );
NOR2_X4 _656_ ( .A1(_270_ ), .A2(_273_ ), .ZN(_274_ ) );
INV_X1 _657_ ( .A(_274_ ), .ZN(_275_ ) );
OAI21_X1 _658_ ( .A(_245_ ), .B1(_275_ ), .B2(_079_ ), .ZN(_276_ ) );
INV_X1 _659_ ( .A(_079_ ), .ZN(_277_ ) );
NOR2_X1 _660_ ( .A1(_274_ ), .A2(_277_ ), .ZN(_278_ ) );
NOR2_X1 _661_ ( .A1(_276_ ), .A2(_278_ ), .ZN(_440_ ) );
NOR2_X4 _662_ ( .A1(_177_ ), .A2(_063_ ), .ZN(_279_ ) );
AND2_X2 _663_ ( .A1(_174_ ), .A2(_030_ ), .ZN(_280_ ) );
OR4_X1 _664_ ( .A1(_279_ ), .A2(_278_ ), .A3(_178_ ), .A4(_280_ ), .ZN(_281_ ) );
OAI22_X1 _665_ ( .A1(_278_ ), .A2(_280_ ), .B1(_279_ ), .B2(_178_ ), .ZN(_282_ ) );
AOI21_X1 _666_ ( .A(_234_ ), .B1(_281_ ), .B2(_282_ ), .ZN(_441_ ) );
NOR4_X1 _667_ ( .A1(_274_ ), .A2(_279_ ), .A3(_178_ ), .A4(_277_ ), .ZN(_283_ ) );
AOI21_X2 _668_ ( .A(_279_ ), .B1(_078_ ), .B2(_280_ ), .ZN(_284_ ) );
INV_X1 _669_ ( .A(_284_ ), .ZN(_285_ ) );
NOR2_X1 _670_ ( .A1(_283_ ), .A2(_285_ ), .ZN(_286_ ) );
INV_X1 _671_ ( .A(_075_ ), .ZN(_287_ ) );
NOR2_X1 _672_ ( .A1(_286_ ), .A2(_287_ ), .ZN(_288_ ) );
NOR3_X1 _673_ ( .A1(_283_ ), .A2(_075_ ), .A3(_285_ ), .ZN(_289_ ) );
NOR3_X1 _674_ ( .A1(_288_ ), .A2(_235_ ), .A3(_289_ ), .ZN(_411_ ) );
NOR2_X4 _675_ ( .A1(_180_ ), .A2(_033_ ), .ZN(_290_ ) );
OR3_X1 _676_ ( .A1(_288_ ), .A2(_290_ ), .A3(_076_ ), .ZN(_291_ ) );
OAI21_X1 _677_ ( .A(_076_ ), .B1(_288_ ), .B2(_290_ ), .ZN(_292_ ) );
AND3_X1 _678_ ( .A1(_291_ ), .A2(_245_ ), .A3(_292_ ), .ZN(_412_ ) );
AND2_X1 _679_ ( .A1(_275_ ), .A2(_080_ ), .ZN(_293_ ) );
NAND2_X2 _680_ ( .A1(_076_ ), .A2(_290_ ), .ZN(_294_ ) );
OAI21_X2 _681_ ( .A(_294_ ), .B1(_181_ ), .B2(_034_ ), .ZN(_295_ ) );
AOI21_X4 _682_ ( .A(_295_ ), .B1(_077_ ), .B2(_285_ ), .ZN(_296_ ) );
INV_X1 _683_ ( .A(_296_ ), .ZN(_297_ ) );
NOR2_X1 _684_ ( .A1(_293_ ), .A2(_297_ ), .ZN(_298_ ) );
INV_X1 _685_ ( .A(_072_ ), .ZN(_299_ ) );
NOR2_X1 _686_ ( .A1(_298_ ), .A2(_299_ ), .ZN(_300_ ) );
AOI211_X4 _687_ ( .A(_072_ ), .B(_297_ ), .C1(_275_ ), .C2(_080_ ), .ZN(_301_ ) );
NOR3_X1 _688_ ( .A1(_300_ ), .A2(_235_ ), .A3(_301_ ), .ZN(_413_ ) );
AND2_X1 _689_ ( .A1(_190_ ), .A2(_003_ ), .ZN(_302_ ) );
OR3_X1 _690_ ( .A1(_300_ ), .A2(_071_ ), .A3(_302_ ), .ZN(_303_ ) );
OAI21_X1 _691_ ( .A(_071_ ), .B1(_300_ ), .B2(_302_ ), .ZN(_304_ ) );
AND3_X1 _692_ ( .A1(_303_ ), .A2(_245_ ), .A3(_304_ ), .ZN(_414_ ) );
INV_X1 _693_ ( .A(_068_ ), .ZN(_305_ ) );
NOR2_X2 _694_ ( .A1(_193_ ), .A2(_036_ ), .ZN(_306_ ) );
NOR4_X1 _695_ ( .A1(_298_ ), .A2(_306_ ), .A3(_194_ ), .A4(_299_ ), .ZN(_307_ ) );
INV_X1 _696_ ( .A(_307_ ), .ZN(_308_ ) );
AOI21_X1 _697_ ( .A(_306_ ), .B1(_071_ ), .B2(_302_ ), .ZN(_309_ ) );
AOI21_X1 _698_ ( .A(_305_ ), .B1(_308_ ), .B2(_309_ ), .ZN(_310_ ) );
AND2_X1 _699_ ( .A1(_308_ ), .A2(_309_ ), .ZN(_311_ ) );
AND2_X1 _700_ ( .A1(_311_ ), .A2(_305_ ), .ZN(_312_ ) );
NOR3_X1 _701_ ( .A1(_310_ ), .A2(_235_ ), .A3(_312_ ), .ZN(_415_ ) );
AND2_X1 _702_ ( .A1(_197_ ), .A2(_005_ ), .ZN(_313_ ) );
OR3_X1 _703_ ( .A1(_310_ ), .A2(_313_ ), .A3(_069_ ), .ZN(_314_ ) );
OAI21_X1 _704_ ( .A(_069_ ), .B1(_310_ ), .B2(_313_ ), .ZN(_315_ ) );
AND3_X1 _705_ ( .A1(_314_ ), .A2(_245_ ), .A3(_315_ ), .ZN(_416_ ) );
NOR2_X4 _706_ ( .A1(_274_ ), .A2(_201_ ), .ZN(_316_ ) );
NOR2_X2 _707_ ( .A1(_296_ ), .A2(_185_ ), .ZN(_317_ ) );
INV_X1 _708_ ( .A(_070_ ), .ZN(_318_ ) );
NOR2_X1 _709_ ( .A1(_318_ ), .A2(_309_ ), .ZN(_319_ ) );
AND2_X1 _710_ ( .A1(_069_ ), .A2(_313_ ), .ZN(_320_ ) );
OR4_X4 _711_ ( .A1(_196_ ), .A2(_317_ ), .A3(_319_ ), .A4(_320_ ), .ZN(_321_ ) );
NOR2_X4 _712_ ( .A1(_316_ ), .A2(_321_ ), .ZN(_322_ ) );
INV_X4 _713_ ( .A(_322_ ), .ZN(_323_ ) );
OAI21_X1 _714_ ( .A(_245_ ), .B1(_323_ ), .B2(_097_ ), .ZN(_324_ ) );
INV_X1 _715_ ( .A(_097_ ), .ZN(_325_ ) );
NOR2_X1 _716_ ( .A1(_322_ ), .A2(_325_ ), .ZN(_326_ ) );
NOR2_X1 _717_ ( .A1(_324_ ), .A2(_326_ ), .ZN(_417_ ) );
AND2_X1 _718_ ( .A1(_140_ ), .A2(_007_ ), .ZN(_327_ ) );
OR4_X1 _719_ ( .A1(_139_ ), .A2(_326_ ), .A3(_138_ ), .A4(_327_ ), .ZN(_328_ ) );
OAI22_X1 _720_ ( .A1(_326_ ), .A2(_327_ ), .B1(_139_ ), .B2(_138_ ), .ZN(_329_ ) );
AOI21_X1 _721_ ( .A(_234_ ), .B1(_328_ ), .B2(_329_ ), .ZN(_418_ ) );
NOR4_X1 _722_ ( .A1(_322_ ), .A2(_139_ ), .A3(_138_ ), .A4(_325_ ), .ZN(_330_ ) );
AOI21_X1 _723_ ( .A(_139_ ), .B1(_096_ ), .B2(_327_ ), .ZN(_331_ ) );
INV_X1 _724_ ( .A(_331_ ), .ZN(_332_ ) );
NOR2_X1 _725_ ( .A1(_330_ ), .A2(_332_ ), .ZN(_333_ ) );
INV_X1 _726_ ( .A(_093_ ), .ZN(_334_ ) );
NOR2_X1 _727_ ( .A1(_333_ ), .A2(_334_ ), .ZN(_335_ ) );
NOR3_X1 _728_ ( .A1(_330_ ), .A2(_093_ ), .A3(_332_ ), .ZN(_336_ ) );
NOR3_X1 _729_ ( .A1(_335_ ), .A2(_235_ ), .A3(_336_ ), .ZN(_419_ ) );
NOR2_X1 _730_ ( .A1(_146_ ), .A2(_041_ ), .ZN(_337_ ) );
OR3_X1 _731_ ( .A1(_335_ ), .A2(_337_ ), .A3(_094_ ), .ZN(_338_ ) );
OAI21_X1 _732_ ( .A(_094_ ), .B1(_335_ ), .B2(_337_ ), .ZN(_339_ ) );
AND3_X1 _733_ ( .A1(_338_ ), .A2(_233_ ), .A3(_339_ ), .ZN(_420_ ) );
AND2_X1 _734_ ( .A1(_323_ ), .A2(_098_ ), .ZN(_340_ ) );
AND2_X1 _735_ ( .A1(_094_ ), .A2(_337_ ), .ZN(_341_ ) );
AOI21_X1 _736_ ( .A(_341_ ), .B1(_010_ ), .B2(_143_ ), .ZN(_342_ ) );
NAND2_X1 _737_ ( .A1(_332_ ), .A2(_095_ ), .ZN(_343_ ) );
AND2_X1 _738_ ( .A1(_342_ ), .A2(_343_ ), .ZN(_344_ ) );
INV_X1 _739_ ( .A(_344_ ), .ZN(_345_ ) );
NOR2_X1 _740_ ( .A1(_340_ ), .A2(_345_ ), .ZN(_346_ ) );
INV_X1 _741_ ( .A(_099_ ), .ZN(_347_ ) );
NOR2_X1 _742_ ( .A1(_346_ ), .A2(_347_ ), .ZN(_348_ ) );
AOI211_X4 _743_ ( .A(_099_ ), .B(_345_ ), .C1(_323_ ), .C2(_098_ ), .ZN(_349_ ) );
NOR3_X1 _744_ ( .A1(_348_ ), .A2(_235_ ), .A3(_349_ ), .ZN(_422_ ) );
AND2_X1 _745_ ( .A1(_134_ ), .A2(_012_ ), .ZN(_350_ ) );
OR3_X1 _746_ ( .A1(_348_ ), .A2(_350_ ), .A3(_100_ ), .ZN(_351_ ) );
OAI21_X1 _747_ ( .A(_100_ ), .B1(_348_ ), .B2(_350_ ), .ZN(_352_ ) );
AND3_X1 _748_ ( .A1(_351_ ), .A2(_233_ ), .A3(_352_ ), .ZN(_423_ ) );
NOR4_X1 _749_ ( .A1(_346_ ), .A2(_133_ ), .A3(_132_ ), .A4(_347_ ), .ZN(_353_ ) );
AOI21_X1 _750_ ( .A(_132_ ), .B1(_100_ ), .B2(_350_ ), .ZN(_354_ ) );
INV_X1 _751_ ( .A(_354_ ), .ZN(_355_ ) );
NOR2_X1 _752_ ( .A1(_353_ ), .A2(_355_ ), .ZN(_356_ ) );
INV_X1 _753_ ( .A(_102_ ), .ZN(_357_ ) );
NOR2_X1 _754_ ( .A1(_356_ ), .A2(_357_ ), .ZN(_358_ ) );
NOR3_X1 _755_ ( .A1(_353_ ), .A2(_102_ ), .A3(_355_ ), .ZN(_359_ ) );
NOR3_X1 _756_ ( .A1(_358_ ), .A2(_235_ ), .A3(_359_ ), .ZN(_424_ ) );
AND2_X1 _757_ ( .A1(_151_ ), .A2(_014_ ), .ZN(_360_ ) );
OR3_X1 _758_ ( .A1(_358_ ), .A2(_360_ ), .A3(_103_ ), .ZN(_361_ ) );
OAI21_X1 _759_ ( .A(_103_ ), .B1(_358_ ), .B2(_360_ ), .ZN(_362_ ) );
AND3_X1 _760_ ( .A1(_361_ ), .A2(_233_ ), .A3(_362_ ), .ZN(_425_ ) );
AND2_X4 _761_ ( .A1(_323_ ), .A2(_106_ ), .ZN(_363_ ) );
AOI21_X1 _762_ ( .A(_149_ ), .B1(_343_ ), .B2(_342_ ), .ZN(_364_ ) );
AND2_X1 _763_ ( .A1(_128_ ), .A2(_015_ ), .ZN(_365_ ) );
AND2_X1 _764_ ( .A1(_355_ ), .A2(_104_ ), .ZN(_366_ ) );
AND2_X1 _765_ ( .A1(_103_ ), .A2(_360_ ), .ZN(_367_ ) );
NOR4_X1 _766_ ( .A1(_364_ ), .A2(_365_ ), .A3(_366_ ), .A4(_367_ ), .ZN(_368_ ) );
INV_X1 _767_ ( .A(_368_ ), .ZN(_369_ ) );
NOR2_X4 _768_ ( .A1(_363_ ), .A2(_369_ ), .ZN(_370_ ) );
INV_X4 _769_ ( .A(_370_ ), .ZN(_371_ ) );
OAI21_X1 _770_ ( .A(_245_ ), .B1(_371_ ), .B2(_117_ ), .ZN(_372_ ) );
INV_X1 _771_ ( .A(_117_ ), .ZN(_373_ ) );
NOR2_X1 _772_ ( .A1(_370_ ), .A2(_373_ ), .ZN(_374_ ) );
NOR2_X1 _773_ ( .A1(_372_ ), .A2(_374_ ), .ZN(_426_ ) );
AND2_X1 _774_ ( .A1(_162_ ), .A2(_016_ ), .ZN(_375_ ) );
OR3_X1 _775_ ( .A1(_374_ ), .A2(_116_ ), .A3(_375_ ), .ZN(_376_ ) );
OAI21_X1 _776_ ( .A(_116_ ), .B1(_374_ ), .B2(_375_ ), .ZN(_377_ ) );
AND3_X1 _777_ ( .A1(_376_ ), .A2(_233_ ), .A3(_377_ ), .ZN(_427_ ) );
INV_X1 _778_ ( .A(_113_ ), .ZN(_378_ ) );
NOR2_X1 _779_ ( .A1(_159_ ), .A2(_049_ ), .ZN(_379_ ) );
NOR4_X1 _780_ ( .A1(_370_ ), .A2(_379_ ), .A3(_160_ ), .A4(_373_ ), .ZN(_380_ ) );
INV_X1 _781_ ( .A(_380_ ), .ZN(_381_ ) );
AOI21_X1 _782_ ( .A(_379_ ), .B1(_116_ ), .B2(_375_ ), .ZN(_382_ ) );
AOI21_X1 _783_ ( .A(_378_ ), .B1(_381_ ), .B2(_382_ ), .ZN(_383_ ) );
AND2_X1 _784_ ( .A1(_381_ ), .A2(_382_ ), .ZN(_384_ ) );
AND2_X1 _785_ ( .A1(_384_ ), .A2(_378_ ), .ZN(_385_ ) );
NOR3_X1 _786_ ( .A1(_383_ ), .A2(_235_ ), .A3(_385_ ), .ZN(_428_ ) );
NOR2_X1 _787_ ( .A1(_168_ ), .A2(_050_ ), .ZN(_386_ ) );
OR3_X1 _788_ ( .A1(_383_ ), .A2(_386_ ), .A3(_114_ ), .ZN(_387_ ) );
OAI21_X1 _789_ ( .A(_114_ ), .B1(_383_ ), .B2(_386_ ), .ZN(_388_ ) );
AND3_X1 _790_ ( .A1(_387_ ), .A2(_233_ ), .A3(_388_ ), .ZN(_429_ ) );
AND2_X4 _791_ ( .A1(_371_ ), .A2(_118_ ), .ZN(_389_ ) );
NAND2_X1 _792_ ( .A1(_114_ ), .A2(_386_ ), .ZN(_390_ ) );
OAI221_X1 _793_ ( .A(_390_ ), .B1(_166_ ), .B2(_051_ ), .C1(_158_ ), .C2(_382_ ), .ZN(_391_ ) );
NOR2_X4 _794_ ( .A1(_389_ ), .A2(_391_ ), .ZN(_392_ ) );
INV_X1 _795_ ( .A(_110_ ), .ZN(_393_ ) );
NOR2_X1 _796_ ( .A1(_392_ ), .A2(_393_ ), .ZN(_394_ ) );
AOI211_X4 _797_ ( .A(_110_ ), .B(_391_ ), .C1(_371_ ), .C2(_118_ ), .ZN(_395_ ) );
NOR3_X1 _798_ ( .A1(_394_ ), .A2(_235_ ), .A3(_395_ ), .ZN(_430_ ) );
NOR2_X1 _799_ ( .A1(_123_ ), .A2(_052_ ), .ZN(_396_ ) );
AND2_X1 _800_ ( .A1(_125_ ), .A2(_021_ ), .ZN(_397_ ) );
OR4_X1 _801_ ( .A1(_396_ ), .A2(_394_ ), .A3(_126_ ), .A4(_397_ ), .ZN(_398_ ) );
OAI22_X1 _802_ ( .A1(_394_ ), .A2(_396_ ), .B1(_126_ ), .B2(_397_ ), .ZN(_399_ ) );
AOI21_X1 _803_ ( .A(_234_ ), .B1(_398_ ), .B2(_399_ ), .ZN(_431_ ) );
INV_X1 _804_ ( .A(_107_ ), .ZN(_400_ ) );
NOR4_X1 _805_ ( .A1(_392_ ), .A2(_393_ ), .A3(_126_ ), .A4(_397_ ), .ZN(_401_ ) );
INV_X1 _806_ ( .A(_401_ ), .ZN(_402_ ) );
AOI21_X1 _807_ ( .A(_397_ ), .B1(_111_ ), .B2(_396_ ), .ZN(_403_ ) );
AOI21_X1 _808_ ( .A(_400_ ), .B1(_402_ ), .B2(_403_ ), .ZN(_404_ ) );
AND2_X1 _809_ ( .A1(_402_ ), .A2(_403_ ), .ZN(_405_ ) );
AND2_X1 _810_ ( .A1(_405_ ), .A2(_400_ ), .ZN(_406_ ) );
NOR3_X1 _811_ ( .A1(_404_ ), .A2(_234_ ), .A3(_406_ ), .ZN(_433_ ) );
NOR2_X1 _812_ ( .A1(_154_ ), .A2(_055_ ), .ZN(_407_ ) );
OR3_X2 _813_ ( .A1(_404_ ), .A2(_407_ ), .A3(_108_ ), .ZN(_408_ ) );
OAI21_X1 _814_ ( .A(_108_ ), .B1(_404_ ), .B2(_407_ ), .ZN(_409_ ) );
AND3_X1 _815_ ( .A1(_408_ ), .A2(_233_ ), .A3(_409_ ), .ZN(_434_ ) );
BUF_X1 _816_ ( .A(\b [0] ), .Z(_032_ ) );
BUF_X1 _817_ ( .A(\a [0] ), .Z(_000_ ) );
BUF_X1 _818_ ( .A(\a [31] ), .Z(_024_ ) );
BUF_X1 _819_ ( .A(\b [31] ), .Z(_056_ ) );
BUF_X1 _820_ ( .A(\a [30] ), .Z(_023_ ) );
BUF_X1 _821_ ( .A(\b [30] ), .Z(_055_ ) );
BUF_X1 _822_ ( .A(\a [29] ), .Z(_021_ ) );
BUF_X1 _823_ ( .A(\b [29] ), .Z(_053_ ) );
BUF_X1 _824_ ( .A(\a [28] ), .Z(_020_ ) );
BUF_X1 _825_ ( .A(\b [28] ), .Z(_052_ ) );
BUF_X1 _826_ ( .A(\a [27] ), .Z(_019_ ) );
BUF_X1 _827_ ( .A(\b [27] ), .Z(_051_ ) );
BUF_X1 _828_ ( .A(\a [26] ), .Z(_018_ ) );
BUF_X1 _829_ ( .A(\b [26] ), .Z(_050_ ) );
BUF_X1 _830_ ( .A(\a [25] ), .Z(_017_ ) );
BUF_X1 _831_ ( .A(\b [25] ), .Z(_049_ ) );
BUF_X1 _832_ ( .A(\a [24] ), .Z(_016_ ) );
BUF_X1 _833_ ( .A(\b [24] ), .Z(_048_ ) );
BUF_X1 _834_ ( .A(\a [23] ), .Z(_015_ ) );
BUF_X1 _835_ ( .A(\b [23] ), .Z(_047_ ) );
BUF_X1 _836_ ( .A(\a [22] ), .Z(_014_ ) );
BUF_X1 _837_ ( .A(\b [22] ), .Z(_046_ ) );
BUF_X1 _838_ ( .A(\a [21] ), .Z(_013_ ) );
BUF_X1 _839_ ( .A(\b [21] ), .Z(_045_ ) );
BUF_X1 _840_ ( .A(\a [20] ), .Z(_012_ ) );
BUF_X1 _841_ ( .A(\b [20] ), .Z(_044_ ) );
BUF_X1 _842_ ( .A(\a [19] ), .Z(_010_ ) );
BUF_X1 _843_ ( .A(\b [19] ), .Z(_042_ ) );
BUF_X1 _844_ ( .A(\a [18] ), .Z(_009_ ) );
BUF_X1 _845_ ( .A(\b [18] ), .Z(_041_ ) );
BUF_X1 _846_ ( .A(\a [17] ), .Z(_008_ ) );
BUF_X1 _847_ ( .A(\b [17] ), .Z(_040_ ) );
BUF_X1 _848_ ( .A(\a [16] ), .Z(_007_ ) );
BUF_X1 _849_ ( .A(\b [16] ), .Z(_039_ ) );
BUF_X1 _850_ ( .A(\a [15] ), .Z(_006_ ) );
BUF_X1 _851_ ( .A(\b [15] ), .Z(_038_ ) );
BUF_X1 _852_ ( .A(\a [14] ), .Z(_005_ ) );
BUF_X1 _853_ ( .A(\b [14] ), .Z(_037_ ) );
BUF_X1 _854_ ( .A(\a [13] ), .Z(_004_ ) );
BUF_X1 _855_ ( .A(\b [13] ), .Z(_036_ ) );
BUF_X1 _856_ ( .A(\a [12] ), .Z(_003_ ) );
BUF_X1 _857_ ( .A(\b [12] ), .Z(_035_ ) );
BUF_X1 _858_ ( .A(\a [11] ), .Z(_002_ ) );
BUF_X1 _859_ ( .A(\b [11] ), .Z(_034_ ) );
BUF_X1 _860_ ( .A(\a [10] ), .Z(_001_ ) );
BUF_X1 _861_ ( .A(\b [10] ), .Z(_033_ ) );
BUF_X1 _862_ ( .A(\a [9] ), .Z(_031_ ) );
BUF_X1 _863_ ( .A(\b [9] ), .Z(_063_ ) );
BUF_X1 _864_ ( .A(\a [8] ), .Z(_030_ ) );
BUF_X1 _865_ ( .A(\b [8] ), .Z(_062_ ) );
BUF_X1 _866_ ( .A(\a [7] ), .Z(_029_ ) );
BUF_X1 _867_ ( .A(\b [7] ), .Z(_061_ ) );
BUF_X1 _868_ ( .A(\a [6] ), .Z(_028_ ) );
BUF_X1 _869_ ( .A(\b [6] ), .Z(_060_ ) );
BUF_X1 _870_ ( .A(\a [5] ), .Z(_027_ ) );
BUF_X1 _871_ ( .A(\b [5] ), .Z(_059_ ) );
BUF_X1 _872_ ( .A(\a [4] ), .Z(_026_ ) );
BUF_X1 _873_ ( .A(\b [4] ), .Z(_058_ ) );
BUF_X1 _874_ ( .A(\a [3] ), .Z(_025_ ) );
BUF_X1 _875_ ( .A(\b [3] ), .Z(_057_ ) );
BUF_X1 _876_ ( .A(\a [2] ), .Z(_022_ ) );
BUF_X1 _877_ ( .A(\b [2] ), .Z(_054_ ) );
BUF_X1 _878_ ( .A(\a [1] ), .Z(_011_ ) );
BUF_X1 _879_ ( .A(\b [1] ), .Z(_043_ ) );
BUF_X1 _880_ ( .A(\ctrl [1] ), .Z(_065_ ) );
BUF_X1 _881_ ( .A(\ctrl [0] ), .Z(_064_ ) );
BUF_X1 _882_ ( .A(\ctrl [2] ), .Z(_066_ ) );
BUF_X1 _883_ ( .A(\ctrl [3] ), .Z(_067_ ) );
BUF_X1 _884_ ( .A(_410_ ), .Z(\result [0] ) );
BUF_X1 _885_ ( .A(_421_ ), .Z(\result [1] ) );
BUF_X1 _886_ ( .A(_432_ ), .Z(\result [2] ) );
BUF_X1 _887_ ( .A(_435_ ), .Z(\result [3] ) );
BUF_X1 _888_ ( .A(_436_ ), .Z(\result [4] ) );
BUF_X1 _889_ ( .A(_437_ ), .Z(\result [5] ) );
BUF_X1 _890_ ( .A(_438_ ), .Z(\result [6] ) );
BUF_X1 _891_ ( .A(_439_ ), .Z(\result [7] ) );
BUF_X1 _892_ ( .A(_440_ ), .Z(\result [8] ) );
BUF_X1 _893_ ( .A(_441_ ), .Z(\result [9] ) );
BUF_X1 _894_ ( .A(_411_ ), .Z(\result [10] ) );
BUF_X1 _895_ ( .A(_412_ ), .Z(\result [11] ) );
BUF_X1 _896_ ( .A(_413_ ), .Z(\result [12] ) );
BUF_X1 _897_ ( .A(_414_ ), .Z(\result [13] ) );
BUF_X1 _898_ ( .A(_415_ ), .Z(\result [14] ) );
BUF_X1 _899_ ( .A(_416_ ), .Z(\result [15] ) );
BUF_X1 _900_ ( .A(_417_ ), .Z(\result [16] ) );
BUF_X1 _901_ ( .A(_418_ ), .Z(\result [17] ) );
BUF_X1 _902_ ( .A(_419_ ), .Z(\result [18] ) );
BUF_X1 _903_ ( .A(_420_ ), .Z(\result [19] ) );
BUF_X1 _904_ ( .A(_422_ ), .Z(\result [20] ) );
BUF_X1 _905_ ( .A(_423_ ), .Z(\result [21] ) );
BUF_X1 _906_ ( .A(_424_ ), .Z(\result [22] ) );
BUF_X1 _907_ ( .A(_425_ ), .Z(\result [23] ) );
BUF_X1 _908_ ( .A(_426_ ), .Z(\result [24] ) );
BUF_X1 _909_ ( .A(_427_ ), .Z(\result [25] ) );
BUF_X1 _910_ ( .A(_428_ ), .Z(\result [26] ) );
BUF_X1 _911_ ( .A(_429_ ), .Z(\result [27] ) );
BUF_X1 _912_ ( .A(_430_ ), .Z(\result [28] ) );
BUF_X1 _913_ ( .A(_431_ ), .Z(\result [29] ) );
BUF_X1 _914_ ( .A(_433_ ), .Z(\result [30] ) );
BUF_X1 _915_ ( .A(_434_ ), .Z(\result [31] ) );

endmodule
