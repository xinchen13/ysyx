module gpio_top_apb(
    input         clock,
    input         reset,
    input  [31:0] in_paddr,
    input         in_psel,
    input         in_penable,
    input  [2:0]  in_pprot,
    input         in_pwrite,
    input  [31:0] in_pwdata,
    input  [3:0]  in_pstrb,
    output        in_pready,
    output [31:0] in_prdata,
    output        in_pslverr,

    output [15:0] gpio_out,
    input  [15:0] gpio_in,
    output [7:0]  gpio_seg_0,
    output [7:0]  gpio_seg_1,
    output [7:0]  gpio_seg_2,
    output [7:0]  gpio_seg_3,
    output [7:0]  gpio_seg_4,
    output [7:0]  gpio_seg_5,
    output [7:0]  gpio_seg_6,
    output [7:0]  gpio_seg_7
);

  assign gpio_out = 16'hf0f0;

endmodule
