module xcore(
    input logic clk,
    input logic rst_n,
);

endmodule
