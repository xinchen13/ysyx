module xcore();
endmodule
