//Generate the verilog at 2024-08-23T20:33:15
module alu0 (
clk,
a,
b,
ctrl,
result
);

input clk ;
input [31:0] a ;
input [31:0] b ;
input [3:0] ctrl ;
output [31:0] result ;

wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire _133_ ;
wire _134_ ;
wire _135_ ;
wire _136_ ;
wire _137_ ;
wire _138_ ;
wire _139_ ;
wire _140_ ;
wire _141_ ;
wire _142_ ;
wire _143_ ;
wire _144_ ;
wire _145_ ;
wire _146_ ;
wire _147_ ;
wire _148_ ;
wire _149_ ;
wire _150_ ;
wire _151_ ;
wire _152_ ;
wire _153_ ;
wire _154_ ;
wire _155_ ;
wire _156_ ;
wire _157_ ;
wire _158_ ;
wire _159_ ;
wire _160_ ;
wire _161_ ;
wire _162_ ;
wire _163_ ;
wire _164_ ;
wire _165_ ;
wire _166_ ;
wire _167_ ;
wire _168_ ;
wire _169_ ;
wire _170_ ;
wire _171_ ;
wire _172_ ;
wire _173_ ;
wire _174_ ;
wire _175_ ;
wire _176_ ;
wire _177_ ;
wire _178_ ;
wire _179_ ;
wire _180_ ;
wire _181_ ;
wire _182_ ;
wire _183_ ;
wire _184_ ;
wire _185_ ;
wire _186_ ;
wire _187_ ;
wire _188_ ;
wire _189_ ;
wire _190_ ;
wire _191_ ;
wire _192_ ;
wire _193_ ;
wire _194_ ;
wire _195_ ;
wire _196_ ;
wire _197_ ;
wire _198_ ;
wire _199_ ;
wire _200_ ;
wire _201_ ;
wire _202_ ;
wire _203_ ;
wire _204_ ;
wire _205_ ;
wire _206_ ;
wire _207_ ;
wire _208_ ;
wire _209_ ;
wire _210_ ;
wire _211_ ;
wire _212_ ;
wire _213_ ;
wire _214_ ;
wire _215_ ;
wire _216_ ;
wire _217_ ;
wire _218_ ;
wire _219_ ;
wire _220_ ;
wire _221_ ;
wire _222_ ;
wire _223_ ;
wire _224_ ;
wire _225_ ;
wire _226_ ;
wire _227_ ;
wire _228_ ;
wire _229_ ;
wire _230_ ;
wire _231_ ;
wire _232_ ;
wire _233_ ;
wire _234_ ;
wire _235_ ;
wire _236_ ;
wire _237_ ;
wire _238_ ;
wire _239_ ;
wire _240_ ;
wire _241_ ;
wire _242_ ;
wire _243_ ;
wire _244_ ;
wire _245_ ;
wire _246_ ;
wire _247_ ;
wire _248_ ;
wire _249_ ;
wire _250_ ;
wire _251_ ;
wire _252_ ;
wire _253_ ;
wire _254_ ;
wire _255_ ;
wire _256_ ;
wire _257_ ;
wire _258_ ;
wire _259_ ;
wire _260_ ;
wire _261_ ;
wire _262_ ;
wire _263_ ;
wire _264_ ;
wire _265_ ;
wire _266_ ;
wire _267_ ;
wire _268_ ;
wire _269_ ;
wire _270_ ;
wire _271_ ;
wire _272_ ;
wire _273_ ;
wire _274_ ;
wire _275_ ;
wire _276_ ;
wire _277_ ;
wire _278_ ;
wire _279_ ;
wire _280_ ;
wire _281_ ;
wire _282_ ;
wire _283_ ;
wire _284_ ;
wire _285_ ;
wire _286_ ;
wire _287_ ;
wire _288_ ;
wire _289_ ;
wire _290_ ;
wire _291_ ;
wire _292_ ;
wire _293_ ;
wire _294_ ;
wire _295_ ;
wire _296_ ;
wire _297_ ;
wire _298_ ;
wire _299_ ;
wire _300_ ;
wire _301_ ;
wire _302_ ;
wire _303_ ;
wire _304_ ;
wire _305_ ;
wire _306_ ;
wire _307_ ;
wire _308_ ;
wire _309_ ;
wire _310_ ;
wire _311_ ;
wire _312_ ;
wire _313_ ;
wire _314_ ;
wire _315_ ;
wire _316_ ;
wire _317_ ;
wire _318_ ;
wire _319_ ;
wire _320_ ;
wire _321_ ;
wire _322_ ;
wire _323_ ;
wire _324_ ;
wire _325_ ;
wire _326_ ;
wire _327_ ;
wire _328_ ;
wire _329_ ;
wire _330_ ;
wire _331_ ;
wire _332_ ;
wire _333_ ;
wire _334_ ;
wire _335_ ;
wire _336_ ;
wire _337_ ;
wire _338_ ;
wire _339_ ;
wire _340_ ;
wire _341_ ;
wire _342_ ;
wire _343_ ;
wire _344_ ;
wire _345_ ;
wire _346_ ;
wire _347_ ;
wire [31:0] a ;
wire [31:0] b ;
wire [3:0] ctrl ;
wire [31:0] result ;


OR3_X1 _348_ ( .A1(_133_ ), .A2(_135_ ), .A3(_136_ ), .ZN(_137_ ) );
AND2_X1 _349_ ( .A1(_130_ ), .A2(_136_ ), .ZN(_138_ ) );
OAI21_X1 _350_ ( .A(_138_ ), .B1(_124_ ), .B2(_128_ ), .ZN(_139_ ) );
AND2_X2 _351_ ( .A1(_136_ ), .A2(_135_ ), .ZN(_140_ ) );
NOR2_X1 _352_ ( .A1(_140_ ), .A2(_073_ ), .ZN(_141_ ) );
AND3_X1 _353_ ( .A1(_137_ ), .A2(_139_ ), .A3(_141_ ), .ZN(_347_ ) );
INV_X1 _354_ ( .A(_063_ ), .ZN(_142_ ) );
AOI21_X2 _355_ ( .A(_140_ ), .B1(_031_ ), .B2(_142_ ), .ZN(_143_ ) );
AND2_X1 _356_ ( .A1(_139_ ), .A2(_143_ ), .ZN(_144_ ) );
INV_X1 _357_ ( .A(_144_ ), .ZN(_145_ ) );
XNOR2_X2 _358_ ( .A(_001_ ), .B(_033_ ), .ZN(_146_ ) );
OAI21_X1 _359_ ( .A(_071_ ), .B1(_145_ ), .B2(_146_ ), .ZN(_147_ ) );
AOI21_X1 _360_ ( .A(_147_ ), .B1(_145_ ), .B2(_146_ ), .ZN(_317_ ) );
INV_X1 _361_ ( .A(_001_ ), .ZN(_148_ ) );
NOR2_X1 _362_ ( .A1(_148_ ), .A2(_033_ ), .ZN(_149_ ) );
AOI21_X1 _363_ ( .A(_149_ ), .B1(_145_ ), .B2(_146_ ), .ZN(_150_ ) );
XNOR2_X2 _364_ ( .A(_002_ ), .B(_034_ ), .ZN(_151_ ) );
XNOR2_X1 _365_ ( .A(_150_ ), .B(_151_ ), .ZN(_152_ ) );
AND3_X1 _366_ ( .A1(_152_ ), .A2(_070_ ), .A3(_069_ ), .ZN(_318_ ) );
AND2_X2 _367_ ( .A1(_151_ ), .A2(_149_ ), .ZN(_153_ ) );
INV_X1 _368_ ( .A(_034_ ), .ZN(_154_ ) );
AOI21_X2 _369_ ( .A(_153_ ), .B1(_002_ ), .B2(_154_ ), .ZN(_155_ ) );
AND2_X1 _370_ ( .A1(_146_ ), .A2(_151_ ), .ZN(_156_ ) );
INV_X1 _371_ ( .A(_156_ ), .ZN(_157_ ) );
OAI21_X1 _372_ ( .A(_155_ ), .B1(_143_ ), .B2(_157_ ), .ZN(_158_ ) );
INV_X4 _373_ ( .A(_129_ ), .ZN(_159_ ) );
AND2_X1 _374_ ( .A1(_138_ ), .A2(_156_ ), .ZN(_160_ ) );
AOI21_X1 _375_ ( .A(_158_ ), .B1(_159_ ), .B2(_160_ ), .ZN(_161_ ) );
XNOR2_X1 _376_ ( .A(_003_ ), .B(_035_ ), .ZN(_162_ ) );
INV_X1 _377_ ( .A(_162_ ), .ZN(_163_ ) );
AND2_X1 _378_ ( .A1(_161_ ), .A2(_163_ ), .ZN(_164_ ) );
NOR2_X2 _379_ ( .A1(_161_ ), .A2(_163_ ), .ZN(_165_ ) );
NOR3_X1 _380_ ( .A1(_164_ ), .A2(_165_ ), .A3(_073_ ), .ZN(_319_ ) );
INV_X1 _381_ ( .A(_003_ ), .ZN(_166_ ) );
NOR2_X1 _382_ ( .A1(_166_ ), .A2(_035_ ), .ZN(_167_ ) );
XNOR2_X2 _383_ ( .A(_004_ ), .B(_036_ ), .ZN(_168_ ) );
NOR3_X1 _384_ ( .A1(_165_ ), .A2(_167_ ), .A3(_168_ ), .ZN(_169_ ) );
AND2_X2 _385_ ( .A1(_165_ ), .A2(_168_ ), .ZN(_170_ ) );
AND2_X2 _386_ ( .A1(_168_ ), .A2(_167_ ), .ZN(_171_ ) );
NOR4_X1 _387_ ( .A1(_169_ ), .A2(_170_ ), .A3(_073_ ), .A4(_171_ ), .ZN(_320_ ) );
INV_X1 _388_ ( .A(_170_ ), .ZN(_172_ ) );
INV_X1 _389_ ( .A(_036_ ), .ZN(_173_ ) );
AOI21_X2 _390_ ( .A(_171_ ), .B1(_004_ ), .B2(_173_ ), .ZN(_174_ ) );
AND2_X2 _391_ ( .A1(_172_ ), .A2(_174_ ), .ZN(_175_ ) );
XNOR2_X1 _392_ ( .A(_005_ ), .B(_037_ ), .ZN(_176_ ) );
INV_X1 _393_ ( .A(_176_ ), .ZN(_177_ ) );
NOR2_X1 _394_ ( .A1(_175_ ), .A2(_177_ ), .ZN(_178_ ) );
INV_X1 _395_ ( .A(_178_ ), .ZN(_179_ ) );
AOI21_X1 _396_ ( .A(_073_ ), .B1(_175_ ), .B2(_177_ ), .ZN(_180_ ) );
AND2_X1 _397_ ( .A1(_179_ ), .A2(_180_ ), .ZN(_321_ ) );
INV_X1 _398_ ( .A(_005_ ), .ZN(_181_ ) );
NOR2_X1 _399_ ( .A1(_181_ ), .A2(_037_ ), .ZN(_182_ ) );
XNOR2_X1 _400_ ( .A(_006_ ), .B(_038_ ), .ZN(_183_ ) );
OR3_X2 _401_ ( .A1(_178_ ), .A2(_182_ ), .A3(_183_ ), .ZN(_184_ ) );
OAI21_X1 _402_ ( .A(_183_ ), .B1(_178_ ), .B2(_182_ ), .ZN(_185_ ) );
AND3_X1 _403_ ( .A1(_184_ ), .A2(_080_ ), .A3(_185_ ), .ZN(_322_ ) );
NAND3_X1 _404_ ( .A1(_168_ ), .A2(_176_ ), .A3(_183_ ), .ZN(_186_ ) );
NOR2_X1 _405_ ( .A1(_186_ ), .A2(_163_ ), .ZN(_187_ ) );
AND3_X4 _406_ ( .A1(_159_ ), .A2(_160_ ), .A3(_187_ ), .ZN(_188_ ) );
AND2_X1 _407_ ( .A1(_158_ ), .A2(_187_ ), .ZN(_189_ ) );
INV_X1 _408_ ( .A(_006_ ), .ZN(_190_ ) );
NOR2_X1 _409_ ( .A1(_190_ ), .A2(_038_ ), .ZN(_191_ ) );
INV_X1 _410_ ( .A(_183_ ), .ZN(_192_ ) );
NOR3_X1 _411_ ( .A1(_174_ ), .A2(_177_ ), .A3(_192_ ), .ZN(_193_ ) );
AND2_X1 _412_ ( .A1(_183_ ), .A2(_182_ ), .ZN(_194_ ) );
NOR4_X1 _413_ ( .A1(_189_ ), .A2(_191_ ), .A3(_193_ ), .A4(_194_ ), .ZN(_195_ ) );
INV_X2 _414_ ( .A(_195_ ), .ZN(_196_ ) );
NOR2_X1 _415_ ( .A1(_188_ ), .A2(_196_ ), .ZN(_197_ ) );
XNOR2_X1 _416_ ( .A(_007_ ), .B(_039_ ), .ZN(_198_ ) );
INV_X1 _417_ ( .A(_198_ ), .ZN(_199_ ) );
NOR2_X1 _418_ ( .A1(_197_ ), .A2(_199_ ), .ZN(_200_ ) );
NOR3_X1 _419_ ( .A1(_188_ ), .A2(_196_ ), .A3(_198_ ), .ZN(_201_ ) );
NOR3_X1 _420_ ( .A1(_200_ ), .A2(_073_ ), .A3(_201_ ), .ZN(_323_ ) );
XNOR2_X1 _421_ ( .A(_008_ ), .B(_040_ ), .ZN(_202_ ) );
NAND2_X1 _422_ ( .A1(_198_ ), .A2(_202_ ), .ZN(_203_ ) );
NOR2_X1 _423_ ( .A1(_197_ ), .A2(_203_ ), .ZN(_204_ ) );
INV_X1 _424_ ( .A(_007_ ), .ZN(_205_ ) );
NOR2_X1 _425_ ( .A1(_205_ ), .A2(_039_ ), .ZN(_206_ ) );
NOR3_X1 _426_ ( .A1(_200_ ), .A2(_206_ ), .A3(_202_ ), .ZN(_207_ ) );
OR2_X1 _427_ ( .A1(_207_ ), .A2(_072_ ), .ZN(_208_ ) );
AOI211_X4 _428_ ( .A(_204_ ), .B(_208_ ), .C1(_206_ ), .C2(_202_ ), .ZN(_324_ ) );
AND2_X1 _429_ ( .A1(_202_ ), .A2(_206_ ), .ZN(_209_ ) );
INV_X1 _430_ ( .A(_040_ ), .ZN(_210_ ) );
AOI21_X1 _431_ ( .A(_209_ ), .B1(_008_ ), .B2(_210_ ), .ZN(_211_ ) );
INV_X1 _432_ ( .A(_211_ ), .ZN(_212_ ) );
NOR2_X1 _433_ ( .A1(_204_ ), .A2(_212_ ), .ZN(_213_ ) );
XNOR2_X1 _434_ ( .A(_009_ ), .B(_041_ ), .ZN(_214_ ) );
INV_X1 _435_ ( .A(_214_ ), .ZN(_215_ ) );
OAI21_X1 _436_ ( .A(_071_ ), .B1(_213_ ), .B2(_215_ ), .ZN(_216_ ) );
AOI21_X1 _437_ ( .A(_216_ ), .B1(_213_ ), .B2(_215_ ), .ZN(_325_ ) );
INV_X1 _438_ ( .A(_009_ ), .ZN(_217_ ) );
NOR2_X1 _439_ ( .A1(_217_ ), .A2(_041_ ), .ZN(_218_ ) );
INV_X1 _440_ ( .A(_218_ ), .ZN(_219_ ) );
OAI21_X1 _441_ ( .A(_219_ ), .B1(_213_ ), .B2(_215_ ), .ZN(_220_ ) );
XNOR2_X1 _442_ ( .A(_010_ ), .B(_042_ ), .ZN(_221_ ) );
OAI21_X1 _443_ ( .A(_071_ ), .B1(_220_ ), .B2(_221_ ), .ZN(_222_ ) );
AOI21_X1 _444_ ( .A(_222_ ), .B1(_220_ ), .B2(_221_ ), .ZN(_326_ ) );
AND2_X1 _445_ ( .A1(_214_ ), .A2(_221_ ), .ZN(_223_ ) );
AND3_X1 _446_ ( .A1(_223_ ), .A2(_198_ ), .A3(_202_ ), .ZN(_224_ ) );
OAI21_X1 _447_ ( .A(_224_ ), .B1(_188_ ), .B2(_196_ ), .ZN(_225_ ) );
NAND2_X1 _448_ ( .A1(_221_ ), .A2(_218_ ), .ZN(_226_ ) );
INV_X1 _449_ ( .A(_010_ ), .ZN(_227_ ) );
OAI21_X1 _450_ ( .A(_226_ ), .B1(_227_ ), .B2(_042_ ), .ZN(_228_ ) );
AOI21_X1 _451_ ( .A(_228_ ), .B1(_212_ ), .B2(_223_ ), .ZN(_229_ ) );
AND2_X2 _452_ ( .A1(_225_ ), .A2(_229_ ), .ZN(_230_ ) );
XNOR2_X1 _453_ ( .A(_012_ ), .B(_044_ ), .ZN(_231_ ) );
INV_X1 _454_ ( .A(_231_ ), .ZN(_232_ ) );
OAI21_X1 _455_ ( .A(_071_ ), .B1(_230_ ), .B2(_232_ ), .ZN(_233_ ) );
AOI21_X1 _456_ ( .A(_233_ ), .B1(_230_ ), .B2(_232_ ), .ZN(_328_ ) );
NOR2_X4 _457_ ( .A1(_230_ ), .A2(_232_ ), .ZN(_234_ ) );
INV_X1 _458_ ( .A(_012_ ), .ZN(_235_ ) );
NOR2_X1 _459_ ( .A1(_235_ ), .A2(_044_ ), .ZN(_236_ ) );
XNOR2_X2 _460_ ( .A(_013_ ), .B(_045_ ), .ZN(_237_ ) );
NOR3_X1 _461_ ( .A1(_234_ ), .A2(_236_ ), .A3(_237_ ), .ZN(_238_ ) );
AND2_X1 _462_ ( .A1(_237_ ), .A2(_236_ ), .ZN(_239_ ) );
OR3_X1 _463_ ( .A1(_238_ ), .A2(_072_ ), .A3(_239_ ), .ZN(_240_ ) );
AOI21_X1 _464_ ( .A(_240_ ), .B1(_234_ ), .B2(_237_ ), .ZN(_329_ ) );
INV_X1 _465_ ( .A(_045_ ), .ZN(_241_ ) );
AOI21_X1 _466_ ( .A(_239_ ), .B1(_013_ ), .B2(_241_ ), .ZN(_242_ ) );
INV_X1 _467_ ( .A(_242_ ), .ZN(_243_ ) );
AOI21_X4 _468_ ( .A(_243_ ), .B1(_234_ ), .B2(_237_ ), .ZN(_244_ ) );
XNOR2_X1 _469_ ( .A(_014_ ), .B(_046_ ), .ZN(_245_ ) );
INV_X1 _470_ ( .A(_245_ ), .ZN(_246_ ) );
NOR2_X2 _471_ ( .A1(_244_ ), .A2(_246_ ), .ZN(_247_ ) );
INV_X1 _472_ ( .A(_247_ ), .ZN(_248_ ) );
AOI21_X1 _473_ ( .A(_073_ ), .B1(_244_ ), .B2(_246_ ), .ZN(_249_ ) );
AND2_X1 _474_ ( .A1(_248_ ), .A2(_249_ ), .ZN(_330_ ) );
INV_X1 _475_ ( .A(_014_ ), .ZN(_250_ ) );
NOR2_X1 _476_ ( .A1(_250_ ), .A2(_046_ ), .ZN(_251_ ) );
XNOR2_X1 _477_ ( .A(_015_ ), .B(_047_ ), .ZN(_252_ ) );
OR3_X4 _478_ ( .A1(_247_ ), .A2(_251_ ), .A3(_252_ ), .ZN(_253_ ) );
OAI21_X1 _479_ ( .A(_252_ ), .B1(_247_ ), .B2(_251_ ), .ZN(_254_ ) );
AND3_X1 _480_ ( .A1(_253_ ), .A2(_080_ ), .A3(_254_ ), .ZN(_331_ ) );
AND2_X1 _481_ ( .A1(_231_ ), .A2(_237_ ), .ZN(_255_ ) );
AND2_X1 _482_ ( .A1(_245_ ), .A2(_252_ ), .ZN(_256_ ) );
AND2_X2 _483_ ( .A1(_255_ ), .A2(_256_ ), .ZN(_257_ ) );
OAI211_X4 _484_ ( .A(_224_ ), .B(_257_ ), .C1(_188_ ), .C2(_196_ ), .ZN(_258_ ) );
NAND2_X1 _485_ ( .A1(_252_ ), .A2(_251_ ), .ZN(_259_ ) );
INV_X1 _486_ ( .A(_015_ ), .ZN(_260_ ) );
INV_X1 _487_ ( .A(_257_ ), .ZN(_261_ ) );
OAI221_X1 _488_ ( .A(_259_ ), .B1(_260_ ), .B2(_047_ ), .C1(_229_ ), .C2(_261_ ), .ZN(_262_ ) );
AOI21_X1 _489_ ( .A(_262_ ), .B1(_243_ ), .B2(_256_ ), .ZN(_263_ ) );
NAND2_X4 _490_ ( .A1(_258_ ), .A2(_263_ ), .ZN(_264_ ) );
XNOR2_X1 _491_ ( .A(_016_ ), .B(_048_ ), .ZN(_265_ ) );
AND2_X1 _492_ ( .A1(_264_ ), .A2(_265_ ), .ZN(_266_ ) );
OAI21_X1 _493_ ( .A(_080_ ), .B1(_264_ ), .B2(_265_ ), .ZN(_267_ ) );
NOR2_X1 _494_ ( .A1(_266_ ), .A2(_267_ ), .ZN(_332_ ) );
XNOR2_X1 _495_ ( .A(_017_ ), .B(_049_ ), .ZN(_268_ ) );
INV_X1 _496_ ( .A(_016_ ), .ZN(_269_ ) );
NOR2_X1 _497_ ( .A1(_269_ ), .A2(_048_ ), .ZN(_270_ ) );
AND2_X1 _498_ ( .A1(_268_ ), .A2(_270_ ), .ZN(_271_ ) );
NOR3_X1 _499_ ( .A1(_266_ ), .A2(_270_ ), .A3(_268_ ), .ZN(_272_ ) );
OR2_X1 _500_ ( .A1(_272_ ), .A2(_072_ ), .ZN(_273_ ) );
AND2_X1 _501_ ( .A1(_265_ ), .A2(_268_ ), .ZN(_274_ ) );
AOI211_X2 _502_ ( .A(_271_ ), .B(_273_ ), .C1(_264_ ), .C2(_274_ ), .ZN(_333_ ) );
INV_X1 _503_ ( .A(_049_ ), .ZN(_275_ ) );
AOI21_X1 _504_ ( .A(_271_ ), .B1(_017_ ), .B2(_275_ ), .ZN(_276_ ) );
INV_X1 _505_ ( .A(_276_ ), .ZN(_277_ ) );
AOI21_X1 _506_ ( .A(_277_ ), .B1(_264_ ), .B2(_274_ ), .ZN(_278_ ) );
XNOR2_X1 _507_ ( .A(_018_ ), .B(_050_ ), .ZN(_279_ ) );
INV_X1 _508_ ( .A(_279_ ), .ZN(_280_ ) );
NOR2_X1 _509_ ( .A1(_278_ ), .A2(_280_ ), .ZN(_281_ ) );
INV_X1 _510_ ( .A(_281_ ), .ZN(_282_ ) );
AOI21_X1 _511_ ( .A(_073_ ), .B1(_278_ ), .B2(_280_ ), .ZN(_283_ ) );
AND2_X1 _512_ ( .A1(_282_ ), .A2(_283_ ), .ZN(_334_ ) );
INV_X1 _513_ ( .A(_018_ ), .ZN(_284_ ) );
NOR2_X1 _514_ ( .A1(_284_ ), .A2(_050_ ), .ZN(_285_ ) );
XNOR2_X1 _515_ ( .A(_019_ ), .B(_051_ ), .ZN(_286_ ) );
OR3_X4 _516_ ( .A1(_281_ ), .A2(_285_ ), .A3(_286_ ), .ZN(_287_ ) );
OAI21_X1 _517_ ( .A(_286_ ), .B1(_281_ ), .B2(_285_ ), .ZN(_288_ ) );
AND3_X1 _518_ ( .A1(_287_ ), .A2(_080_ ), .A3(_288_ ), .ZN(_335_ ) );
AND2_X1 _519_ ( .A1(_279_ ), .A2(_286_ ), .ZN(_289_ ) );
NAND3_X4 _520_ ( .A1(_264_ ), .A2(_274_ ), .A3(_289_ ), .ZN(_290_ ) );
AND2_X1 _521_ ( .A1(_286_ ), .A2(_285_ ), .ZN(_291_ ) );
INV_X1 _522_ ( .A(_051_ ), .ZN(_292_ ) );
AOI221_X4 _523_ ( .A(_291_ ), .B1(_019_ ), .B2(_292_ ), .C1(_277_ ), .C2(_289_ ), .ZN(_293_ ) );
AND2_X4 _524_ ( .A1(_290_ ), .A2(_293_ ), .ZN(_294_ ) );
XNOR2_X1 _525_ ( .A(_020_ ), .B(_052_ ), .ZN(_295_ ) );
INV_X1 _526_ ( .A(_295_ ), .ZN(_296_ ) );
NOR2_X2 _527_ ( .A1(_294_ ), .A2(_296_ ), .ZN(_297_ ) );
AND3_X1 _528_ ( .A1(_290_ ), .A2(_293_ ), .A3(_296_ ), .ZN(_298_ ) );
NOR3_X1 _529_ ( .A1(_297_ ), .A2(_073_ ), .A3(_298_ ), .ZN(_336_ ) );
INV_X1 _530_ ( .A(_020_ ), .ZN(_299_ ) );
NOR2_X1 _531_ ( .A1(_299_ ), .A2(_052_ ), .ZN(_300_ ) );
XNOR2_X1 _532_ ( .A(_021_ ), .B(_053_ ), .ZN(_301_ ) );
OR3_X4 _533_ ( .A1(_297_ ), .A2(_300_ ), .A3(_301_ ), .ZN(_302_ ) );
NAND2_X1 _534_ ( .A1(_295_ ), .A2(_301_ ), .ZN(_303_ ) );
OR2_X4 _535_ ( .A1(_294_ ), .A2(_303_ ), .ZN(_304_ ) );
NAND2_X1 _536_ ( .A1(_301_ ), .A2(_300_ ), .ZN(_305_ ) );
AND4_X1 _537_ ( .A1(_080_ ), .A2(_302_ ), .A3(_304_ ), .A4(_305_ ), .ZN(_337_ ) );
INV_X1 _538_ ( .A(_053_ ), .ZN(_306_ ) );
NAND2_X1 _539_ ( .A1(_306_ ), .A2(_021_ ), .ZN(_307_ ) );
AND3_X4 _540_ ( .A1(_304_ ), .A2(_307_ ), .A3(_305_ ), .ZN(_308_ ) );
XOR2_X1 _541_ ( .A(_023_ ), .B(_055_ ), .Z(_309_ ) );
OAI21_X1 _542_ ( .A(_071_ ), .B1(_308_ ), .B2(_309_ ), .ZN(_310_ ) );
AOI21_X1 _543_ ( .A(_310_ ), .B1(_308_ ), .B2(_309_ ), .ZN(_339_ ) );
INV_X1 _544_ ( .A(_055_ ), .ZN(_311_ ) );
NAND2_X1 _545_ ( .A1(_311_ ), .A2(_023_ ), .ZN(_312_ ) );
OAI21_X4 _546_ ( .A(_312_ ), .B1(_308_ ), .B2(_309_ ), .ZN(_313_ ) );
XNOR2_X1 _547_ ( .A(_024_ ), .B(_056_ ), .ZN(_314_ ) );
OAI21_X1 _548_ ( .A(_071_ ), .B1(_313_ ), .B2(_314_ ), .ZN(_315_ ) );
AOI21_X1 _549_ ( .A(_315_ ), .B1(_313_ ), .B2(_314_ ), .ZN(_340_ ) );
INV_X1 _550_ ( .A(_067_ ), .ZN(_068_ ) );
NOR2_X1 _551_ ( .A1(_068_ ), .A2(_066_ ), .ZN(_069_ ) );
NOR2_X1 _552_ ( .A1(_065_ ), .A2(_064_ ), .ZN(_070_ ) );
AND2_X2 _553_ ( .A1(_069_ ), .A2(_070_ ), .ZN(_071_ ) );
INV_X1 _554_ ( .A(_071_ ), .ZN(_072_ ) );
BUF_X4 _555_ ( .A(_072_ ), .Z(_073_ ) );
INV_X1 _556_ ( .A(_000_ ), .ZN(_074_ ) );
NAND2_X2 _557_ ( .A1(_074_ ), .A2(_032_ ), .ZN(_075_ ) );
OR2_X1 _558_ ( .A1(_074_ ), .A2(_032_ ), .ZN(_076_ ) );
AOI21_X1 _559_ ( .A(_073_ ), .B1(_075_ ), .B2(_076_ ), .ZN(_316_ ) );
XNOR2_X2 _560_ ( .A(_011_ ), .B(_043_ ), .ZN(_077_ ) );
OAI211_X2 _561_ ( .A(_070_ ), .B(_069_ ), .C1(_077_ ), .C2(_075_ ), .ZN(_078_ ) );
AND2_X4 _562_ ( .A1(_077_ ), .A2(_075_ ), .ZN(_079_ ) );
NOR2_X1 _563_ ( .A1(_078_ ), .A2(_079_ ), .ZN(_327_ ) );
BUF_X2 _564_ ( .A(_071_ ), .Z(_080_ ) );
INV_X1 _565_ ( .A(_043_ ), .ZN(_081_ ) );
AOI21_X4 _566_ ( .A(_079_ ), .B1(_011_ ), .B2(_081_ ), .ZN(_082_ ) );
XNOR2_X1 _567_ ( .A(_022_ ), .B(_054_ ), .ZN(_083_ ) );
INV_X1 _568_ ( .A(_083_ ), .ZN(_084_ ) );
OAI21_X1 _569_ ( .A(_080_ ), .B1(_082_ ), .B2(_084_ ), .ZN(_085_ ) );
AOI21_X1 _570_ ( .A(_085_ ), .B1(_082_ ), .B2(_084_ ), .ZN(_338_ ) );
NOR2_X1 _571_ ( .A1(_082_ ), .A2(_084_ ), .ZN(_086_ ) );
INV_X1 _572_ ( .A(_022_ ), .ZN(_087_ ) );
NOR2_X2 _573_ ( .A1(_087_ ), .A2(_054_ ), .ZN(_088_ ) );
XNOR2_X2 _574_ ( .A(_025_ ), .B(_057_ ), .ZN(_089_ ) );
NOR3_X1 _575_ ( .A1(_086_ ), .A2(_088_ ), .A3(_089_ ), .ZN(_090_ ) );
NAND2_X1 _576_ ( .A1(_083_ ), .A2(_089_ ), .ZN(_091_ ) );
NOR2_X4 _577_ ( .A1(_082_ ), .A2(_091_ ), .ZN(_092_ ) );
AND2_X4 _578_ ( .A1(_089_ ), .A2(_088_ ), .ZN(_093_ ) );
NOR4_X1 _579_ ( .A1(_090_ ), .A2(_073_ ), .A3(_092_ ), .A4(_093_ ), .ZN(_341_ ) );
INV_X1 _580_ ( .A(_057_ ), .ZN(_094_ ) );
AOI21_X2 _581_ ( .A(_093_ ), .B1(_025_ ), .B2(_094_ ), .ZN(_095_ ) );
INV_X2 _582_ ( .A(_095_ ), .ZN(_096_ ) );
NOR2_X4 _583_ ( .A1(_092_ ), .A2(_096_ ), .ZN(_097_ ) );
INV_X4 _584_ ( .A(_097_ ), .ZN(_098_ ) );
XNOR2_X1 _585_ ( .A(_026_ ), .B(_058_ ), .ZN(_099_ ) );
OAI21_X1 _586_ ( .A(_080_ ), .B1(_098_ ), .B2(_099_ ), .ZN(_100_ ) );
INV_X1 _587_ ( .A(_099_ ), .ZN(_101_ ) );
NOR2_X1 _588_ ( .A1(_097_ ), .A2(_101_ ), .ZN(_102_ ) );
NOR2_X1 _589_ ( .A1(_100_ ), .A2(_102_ ), .ZN(_342_ ) );
INV_X1 _590_ ( .A(_026_ ), .ZN(_103_ ) );
NOR2_X2 _591_ ( .A1(_103_ ), .A2(_058_ ), .ZN(_104_ ) );
XNOR2_X2 _592_ ( .A(_027_ ), .B(_059_ ), .ZN(_105_ ) );
OR3_X1 _593_ ( .A1(_102_ ), .A2(_104_ ), .A3(_105_ ), .ZN(_106_ ) );
AND2_X4 _594_ ( .A1(_105_ ), .A2(_104_ ), .ZN(_107_ ) );
AND2_X1 _595_ ( .A1(_099_ ), .A2(_105_ ), .ZN(_108_ ) );
AOI211_X4 _596_ ( .A(_072_ ), .B(_107_ ), .C1(_098_ ), .C2(_108_ ), .ZN(_109_ ) );
AND2_X1 _597_ ( .A1(_106_ ), .A2(_109_ ), .ZN(_343_ ) );
INV_X1 _598_ ( .A(_059_ ), .ZN(_110_ ) );
AOI21_X4 _599_ ( .A(_107_ ), .B1(_027_ ), .B2(_110_ ), .ZN(_111_ ) );
INV_X2 _600_ ( .A(_111_ ), .ZN(_112_ ) );
AOI21_X1 _601_ ( .A(_112_ ), .B1(_098_ ), .B2(_108_ ), .ZN(_113_ ) );
XNOR2_X1 _602_ ( .A(_028_ ), .B(_060_ ), .ZN(_114_ ) );
INV_X1 _603_ ( .A(_114_ ), .ZN(_115_ ) );
OAI21_X1 _604_ ( .A(_080_ ), .B1(_113_ ), .B2(_115_ ), .ZN(_116_ ) );
AOI21_X1 _605_ ( .A(_116_ ), .B1(_113_ ), .B2(_115_ ), .ZN(_344_ ) );
NOR2_X1 _606_ ( .A1(_113_ ), .A2(_115_ ), .ZN(_117_ ) );
INV_X1 _607_ ( .A(_028_ ), .ZN(_118_ ) );
NOR2_X1 _608_ ( .A1(_118_ ), .A2(_060_ ), .ZN(_119_ ) );
OR2_X1 _609_ ( .A1(_117_ ), .A2(_119_ ), .ZN(_120_ ) );
XNOR2_X2 _610_ ( .A(_029_ ), .B(_061_ ), .ZN(_121_ ) );
OAI21_X1 _611_ ( .A(_080_ ), .B1(_120_ ), .B2(_121_ ), .ZN(_122_ ) );
AOI21_X1 _612_ ( .A(_122_ ), .B1(_120_ ), .B2(_121_ ), .ZN(_345_ ) );
AND2_X1 _613_ ( .A1(_114_ ), .A2(_121_ ), .ZN(_123_ ) );
AND3_X4 _614_ ( .A1(_098_ ), .A2(_108_ ), .A3(_123_ ), .ZN(_124_ ) );
AND2_X1 _615_ ( .A1(_121_ ), .A2(_119_ ), .ZN(_125_ ) );
INV_X1 _616_ ( .A(_061_ ), .ZN(_126_ ) );
AOI221_X1 _617_ ( .A(_125_ ), .B1(_029_ ), .B2(_126_ ), .C1(_112_ ), .C2(_123_ ), .ZN(_127_ ) );
INV_X1 _618_ ( .A(_127_ ), .ZN(_128_ ) );
NOR2_X4 _619_ ( .A1(_124_ ), .A2(_128_ ), .ZN(_129_ ) );
XNOR2_X1 _620_ ( .A(_030_ ), .B(_062_ ), .ZN(_130_ ) );
INV_X1 _621_ ( .A(_130_ ), .ZN(_131_ ) );
OAI21_X1 _622_ ( .A(_080_ ), .B1(_129_ ), .B2(_131_ ), .ZN(_132_ ) );
AOI21_X1 _623_ ( .A(_132_ ), .B1(_129_ ), .B2(_131_ ), .ZN(_346_ ) );
NOR2_X1 _624_ ( .A1(_129_ ), .A2(_131_ ), .ZN(_133_ ) );
INV_X1 _625_ ( .A(_030_ ), .ZN(_134_ ) );
NOR2_X1 _626_ ( .A1(_134_ ), .A2(_062_ ), .ZN(_135_ ) );
XNOR2_X2 _627_ ( .A(_031_ ), .B(_063_ ), .ZN(_136_ ) );
BUF_X1 _628_ ( .A(\a [0] ), .Z(_000_ ) );
BUF_X1 _629_ ( .A(\b [0] ), .Z(_032_ ) );
BUF_X1 _630_ ( .A(\ctrl [1] ), .Z(_065_ ) );
BUF_X1 _631_ ( .A(\ctrl [0] ), .Z(_064_ ) );
BUF_X1 _632_ ( .A(\ctrl [2] ), .Z(_066_ ) );
BUF_X1 _633_ ( .A(\ctrl [3] ), .Z(_067_ ) );
BUF_X1 _634_ ( .A(_316_ ), .Z(\result [0] ) );
BUF_X1 _635_ ( .A(\a [1] ), .Z(_011_ ) );
BUF_X1 _636_ ( .A(\b [1] ), .Z(_043_ ) );
BUF_X1 _637_ ( .A(_327_ ), .Z(\result [1] ) );
BUF_X1 _638_ ( .A(\a [2] ), .Z(_022_ ) );
BUF_X1 _639_ ( .A(\b [2] ), .Z(_054_ ) );
BUF_X1 _640_ ( .A(_338_ ), .Z(\result [2] ) );
BUF_X1 _641_ ( .A(\a [3] ), .Z(_025_ ) );
BUF_X1 _642_ ( .A(\b [3] ), .Z(_057_ ) );
BUF_X1 _643_ ( .A(_341_ ), .Z(\result [3] ) );
BUF_X1 _644_ ( .A(\a [4] ), .Z(_026_ ) );
BUF_X1 _645_ ( .A(\b [4] ), .Z(_058_ ) );
BUF_X1 _646_ ( .A(_342_ ), .Z(\result [4] ) );
BUF_X1 _647_ ( .A(\a [5] ), .Z(_027_ ) );
BUF_X1 _648_ ( .A(\b [5] ), .Z(_059_ ) );
BUF_X1 _649_ ( .A(_343_ ), .Z(\result [5] ) );
BUF_X1 _650_ ( .A(\a [6] ), .Z(_028_ ) );
BUF_X1 _651_ ( .A(\b [6] ), .Z(_060_ ) );
BUF_X1 _652_ ( .A(_344_ ), .Z(\result [6] ) );
BUF_X1 _653_ ( .A(\a [7] ), .Z(_029_ ) );
BUF_X1 _654_ ( .A(\b [7] ), .Z(_061_ ) );
BUF_X1 _655_ ( .A(_345_ ), .Z(\result [7] ) );
BUF_X1 _656_ ( .A(\a [8] ), .Z(_030_ ) );
BUF_X1 _657_ ( .A(\b [8] ), .Z(_062_ ) );
BUF_X1 _658_ ( .A(_346_ ), .Z(\result [8] ) );
BUF_X1 _659_ ( .A(\a [9] ), .Z(_031_ ) );
BUF_X1 _660_ ( .A(\b [9] ), .Z(_063_ ) );
BUF_X1 _661_ ( .A(_347_ ), .Z(\result [9] ) );
BUF_X1 _662_ ( .A(\a [10] ), .Z(_001_ ) );
BUF_X1 _663_ ( .A(\b [10] ), .Z(_033_ ) );
BUF_X1 _664_ ( .A(_317_ ), .Z(\result [10] ) );
BUF_X1 _665_ ( .A(\a [11] ), .Z(_002_ ) );
BUF_X1 _666_ ( .A(\b [11] ), .Z(_034_ ) );
BUF_X1 _667_ ( .A(_318_ ), .Z(\result [11] ) );
BUF_X1 _668_ ( .A(\a [12] ), .Z(_003_ ) );
BUF_X1 _669_ ( .A(\b [12] ), .Z(_035_ ) );
BUF_X1 _670_ ( .A(_319_ ), .Z(\result [12] ) );
BUF_X1 _671_ ( .A(\a [13] ), .Z(_004_ ) );
BUF_X1 _672_ ( .A(\b [13] ), .Z(_036_ ) );
BUF_X1 _673_ ( .A(_320_ ), .Z(\result [13] ) );
BUF_X1 _674_ ( .A(\a [14] ), .Z(_005_ ) );
BUF_X1 _675_ ( .A(\b [14] ), .Z(_037_ ) );
BUF_X1 _676_ ( .A(_321_ ), .Z(\result [14] ) );
BUF_X1 _677_ ( .A(\a [15] ), .Z(_006_ ) );
BUF_X1 _678_ ( .A(\b [15] ), .Z(_038_ ) );
BUF_X1 _679_ ( .A(_322_ ), .Z(\result [15] ) );
BUF_X1 _680_ ( .A(\a [16] ), .Z(_007_ ) );
BUF_X1 _681_ ( .A(\b [16] ), .Z(_039_ ) );
BUF_X1 _682_ ( .A(_323_ ), .Z(\result [16] ) );
BUF_X1 _683_ ( .A(\a [17] ), .Z(_008_ ) );
BUF_X1 _684_ ( .A(\b [17] ), .Z(_040_ ) );
BUF_X1 _685_ ( .A(_324_ ), .Z(\result [17] ) );
BUF_X1 _686_ ( .A(\a [18] ), .Z(_009_ ) );
BUF_X1 _687_ ( .A(\b [18] ), .Z(_041_ ) );
BUF_X1 _688_ ( .A(_325_ ), .Z(\result [18] ) );
BUF_X1 _689_ ( .A(\a [19] ), .Z(_010_ ) );
BUF_X1 _690_ ( .A(\b [19] ), .Z(_042_ ) );
BUF_X1 _691_ ( .A(_326_ ), .Z(\result [19] ) );
BUF_X1 _692_ ( .A(\a [20] ), .Z(_012_ ) );
BUF_X1 _693_ ( .A(\b [20] ), .Z(_044_ ) );
BUF_X1 _694_ ( .A(_328_ ), .Z(\result [20] ) );
BUF_X1 _695_ ( .A(\a [21] ), .Z(_013_ ) );
BUF_X1 _696_ ( .A(\b [21] ), .Z(_045_ ) );
BUF_X1 _697_ ( .A(_329_ ), .Z(\result [21] ) );
BUF_X1 _698_ ( .A(\a [22] ), .Z(_014_ ) );
BUF_X1 _699_ ( .A(\b [22] ), .Z(_046_ ) );
BUF_X1 _700_ ( .A(_330_ ), .Z(\result [22] ) );
BUF_X1 _701_ ( .A(\a [23] ), .Z(_015_ ) );
BUF_X1 _702_ ( .A(\b [23] ), .Z(_047_ ) );
BUF_X1 _703_ ( .A(_331_ ), .Z(\result [23] ) );
BUF_X1 _704_ ( .A(\a [24] ), .Z(_016_ ) );
BUF_X1 _705_ ( .A(\b [24] ), .Z(_048_ ) );
BUF_X1 _706_ ( .A(_332_ ), .Z(\result [24] ) );
BUF_X1 _707_ ( .A(\a [25] ), .Z(_017_ ) );
BUF_X1 _708_ ( .A(\b [25] ), .Z(_049_ ) );
BUF_X1 _709_ ( .A(_333_ ), .Z(\result [25] ) );
BUF_X1 _710_ ( .A(\a [26] ), .Z(_018_ ) );
BUF_X1 _711_ ( .A(\b [26] ), .Z(_050_ ) );
BUF_X1 _712_ ( .A(_334_ ), .Z(\result [26] ) );
BUF_X1 _713_ ( .A(\a [27] ), .Z(_019_ ) );
BUF_X1 _714_ ( .A(\b [27] ), .Z(_051_ ) );
BUF_X1 _715_ ( .A(_335_ ), .Z(\result [27] ) );
BUF_X1 _716_ ( .A(\a [28] ), .Z(_020_ ) );
BUF_X1 _717_ ( .A(\b [28] ), .Z(_052_ ) );
BUF_X1 _718_ ( .A(_336_ ), .Z(\result [28] ) );
BUF_X1 _719_ ( .A(\a [29] ), .Z(_021_ ) );
BUF_X1 _720_ ( .A(\b [29] ), .Z(_053_ ) );
BUF_X1 _721_ ( .A(_337_ ), .Z(\result [29] ) );
BUF_X1 _722_ ( .A(\a [30] ), .Z(_023_ ) );
BUF_X1 _723_ ( .A(\b [30] ), .Z(_055_ ) );
BUF_X1 _724_ ( .A(_339_ ), .Z(\result [30] ) );
BUF_X1 _725_ ( .A(\a [31] ), .Z(_024_ ) );
BUF_X1 _726_ ( .A(\b [31] ), .Z(_056_ ) );
BUF_X1 _727_ ( .A(_340_ ), .Z(\result [31] ) );

endmodule
