//Generate the verilog at 2024-07-13T10:24:20
module top (
clk,
overflow,
ps2_clk,
ps2_data,
rst_n,
ascii_seg,
count_seg,
scan_code_seg
);

input clk ;
output overflow ;
input ps2_clk ;
input ps2_data ;
input rst_n ;
output [15:0] ascii_seg ;
output [15:0] count_seg ;
output [15:0] scan_code_seg ;

wire _000_ ;
wire _001_ ;
wire _002_ ;
wire _003_ ;
wire _004_ ;
wire _005_ ;
wire _006_ ;
wire _007_ ;
wire _008_ ;
wire _009_ ;
wire _010_ ;
wire _011_ ;
wire _012_ ;
wire _013_ ;
wire _014_ ;
wire _015_ ;
wire _016_ ;
wire _017_ ;
wire _018_ ;
wire _019_ ;
wire _020_ ;
wire _021_ ;
wire _022_ ;
wire _023_ ;
wire _024_ ;
wire _025_ ;
wire _026_ ;
wire _027_ ;
wire _028_ ;
wire _029_ ;
wire _030_ ;
wire _031_ ;
wire _032_ ;
wire _033_ ;
wire _034_ ;
wire _035_ ;
wire _036_ ;
wire _037_ ;
wire _038_ ;
wire _039_ ;
wire _040_ ;
wire _041_ ;
wire _042_ ;
wire _043_ ;
wire _044_ ;
wire _045_ ;
wire _046_ ;
wire _047_ ;
wire _048_ ;
wire _049_ ;
wire _050_ ;
wire _051_ ;
wire _052_ ;
wire _053_ ;
wire _054_ ;
wire _055_ ;
wire _056_ ;
wire _057_ ;
wire _058_ ;
wire _059_ ;
wire _060_ ;
wire _061_ ;
wire _062_ ;
wire _063_ ;
wire _064_ ;
wire _065_ ;
wire _066_ ;
wire _067_ ;
wire _068_ ;
wire _069_ ;
wire _070_ ;
wire _071_ ;
wire _072_ ;
wire _073_ ;
wire _074_ ;
wire _075_ ;
wire _076_ ;
wire _077_ ;
wire _078_ ;
wire _079_ ;
wire _080_ ;
wire _081_ ;
wire _082_ ;
wire _083_ ;
wire _084_ ;
wire _085_ ;
wire _086_ ;
wire _087_ ;
wire _088_ ;
wire _089_ ;
wire _090_ ;
wire _091_ ;
wire _092_ ;
wire _093_ ;
wire _094_ ;
wire _095_ ;
wire _096_ ;
wire _097_ ;
wire _098_ ;
wire _099_ ;
wire _100_ ;
wire _101_ ;
wire _102_ ;
wire _103_ ;
wire _104_ ;
wire _105_ ;
wire _106_ ;
wire _107_ ;
wire _108_ ;
wire _109_ ;
wire _110_ ;
wire _111_ ;
wire _112_ ;
wire _113_ ;
wire _114_ ;
wire _115_ ;
wire _116_ ;
wire _117_ ;
wire _118_ ;
wire _119_ ;
wire _120_ ;
wire _121_ ;
wire _122_ ;
wire _123_ ;
wire _124_ ;
wire _125_ ;
wire _126_ ;
wire _127_ ;
wire _128_ ;
wire _129_ ;
wire _130_ ;
wire _131_ ;
wire _132_ ;
wire _133_ ;
wire _134_ ;
wire _135_ ;
wire _136_ ;
wire _137_ ;
wire _138_ ;
wire _139_ ;
wire _140_ ;
wire _141_ ;
wire _142_ ;
wire count_en ;
wire display_en ;
wire ready ;
wire \u_ascii_h/_00_ ;
wire \u_ascii_h/_01_ ;
wire \u_ascii_h/_02_ ;
wire \u_ascii_h/_03_ ;
wire \u_ascii_h/_04_ ;
wire \u_ascii_h/_05_ ;
wire \u_ascii_h/_06_ ;
wire \u_ascii_h/_07_ ;
wire \u_ascii_h/_08_ ;
wire \u_ascii_h/_09_ ;
wire \u_ascii_h/_10_ ;
wire \u_ascii_h/_11_ ;
wire \u_ascii_h/_12_ ;
wire \u_ascii_h/_13_ ;
wire \u_ascii_h/_14_ ;
wire \u_ascii_h/_15_ ;
wire \u_ascii_h/_16_ ;
wire \u_ascii_h/_17_ ;
wire \u_ascii_h/_18_ ;
wire \u_ascii_h/_19_ ;
wire \u_ascii_h/_20_ ;
wire \u_ascii_h/_21_ ;
wire \u_ascii_h/_22_ ;
wire \u_ascii_h/_23_ ;
wire \u_ascii_h/_24_ ;
wire \u_ascii_h/_25_ ;
wire \u_ascii_h/_26_ ;
wire \u_ascii_h/_27_ ;
wire \u_ascii_h/_28_ ;
wire \u_ascii_h/_29_ ;
wire \u_ascii_h/_30_ ;
wire \u_ascii_h/_31_ ;
wire \u_ascii_h/_32_ ;
wire \u_ascii_h/_33_ ;
wire \u_ascii_h/_34_ ;
wire \u_ascii_h/_35_ ;
wire \u_ascii_h/_36_ ;
wire \u_ascii_h/_37_ ;
wire \u_ascii_h/_38_ ;
wire \u_ascii_h/_39_ ;
wire \u_ascii_h/_40_ ;
wire \u_ascii_h/_41_ ;
wire \u_ascii_h/_42_ ;
wire \u_ascii_l/_00_ ;
wire \u_ascii_l/_01_ ;
wire \u_ascii_l/_02_ ;
wire \u_ascii_l/_03_ ;
wire \u_ascii_l/_04_ ;
wire \u_ascii_l/_05_ ;
wire \u_ascii_l/_06_ ;
wire \u_ascii_l/_07_ ;
wire \u_ascii_l/_08_ ;
wire \u_ascii_l/_09_ ;
wire \u_ascii_l/_10_ ;
wire \u_ascii_l/_11_ ;
wire \u_ascii_l/_12_ ;
wire \u_ascii_l/_13_ ;
wire \u_ascii_l/_14_ ;
wire \u_ascii_l/_15_ ;
wire \u_ascii_l/_16_ ;
wire \u_ascii_l/_17_ ;
wire \u_ascii_l/_18_ ;
wire \u_ascii_l/_19_ ;
wire \u_ascii_l/_20_ ;
wire \u_ascii_l/_21_ ;
wire \u_ascii_l/_22_ ;
wire \u_ascii_l/_23_ ;
wire \u_ascii_l/_24_ ;
wire \u_ascii_l/_25_ ;
wire \u_ascii_l/_26_ ;
wire \u_ascii_l/_27_ ;
wire \u_ascii_l/_28_ ;
wire \u_ascii_l/_29_ ;
wire \u_ascii_l/_30_ ;
wire \u_ascii_l/_31_ ;
wire \u_ascii_l/_32_ ;
wire \u_ascii_l/_33_ ;
wire \u_ascii_l/_34_ ;
wire \u_ascii_l/_35_ ;
wire \u_ascii_l/_36_ ;
wire \u_ascii_l/_37_ ;
wire \u_ascii_l/_38_ ;
wire \u_ascii_l/_39_ ;
wire \u_ascii_l/_40_ ;
wire \u_ascii_l/_41_ ;
wire \u_ascii_l/_42_ ;
wire \u_count_h/_00_ ;
wire \u_count_h/_01_ ;
wire \u_count_h/_02_ ;
wire \u_count_h/_03_ ;
wire \u_count_h/_04_ ;
wire \u_count_h/_05_ ;
wire \u_count_h/_06_ ;
wire \u_count_h/_07_ ;
wire \u_count_h/_08_ ;
wire \u_count_h/_09_ ;
wire \u_count_h/_10_ ;
wire \u_count_h/_11_ ;
wire \u_count_h/_12_ ;
wire \u_count_h/_13_ ;
wire \u_count_h/_14_ ;
wire \u_count_h/_15_ ;
wire \u_count_h/_16_ ;
wire \u_count_h/_17_ ;
wire \u_count_h/_18_ ;
wire \u_count_h/_19_ ;
wire \u_count_h/_20_ ;
wire \u_count_h/_21_ ;
wire \u_count_h/_22_ ;
wire \u_count_h/_23_ ;
wire \u_count_h/_24_ ;
wire \u_count_h/_25_ ;
wire \u_count_h/_26_ ;
wire \u_count_h/_27_ ;
wire \u_count_h/_28_ ;
wire \u_count_h/_29_ ;
wire \u_count_h/_30_ ;
wire \u_count_h/_31_ ;
wire \u_count_h/_32_ ;
wire \u_count_h/_33_ ;
wire \u_count_h/_34_ ;
wire \u_count_h/_35_ ;
wire \u_count_h/_36_ ;
wire \u_count_h/_37_ ;
wire \u_count_h/_38_ ;
wire \u_count_h/_39_ ;
wire \u_count_h/_40_ ;
wire \u_count_h/_41_ ;
wire \u_count_h/_42_ ;
wire \u_count_l/_00_ ;
wire \u_count_l/_01_ ;
wire \u_count_l/_02_ ;
wire \u_count_l/_03_ ;
wire \u_count_l/_04_ ;
wire \u_count_l/_05_ ;
wire \u_count_l/_06_ ;
wire \u_count_l/_07_ ;
wire \u_count_l/_08_ ;
wire \u_count_l/_09_ ;
wire \u_count_l/_10_ ;
wire \u_count_l/_11_ ;
wire \u_count_l/_12_ ;
wire \u_count_l/_13_ ;
wire \u_count_l/_14_ ;
wire \u_count_l/_15_ ;
wire \u_count_l/_16_ ;
wire \u_count_l/_17_ ;
wire \u_count_l/_18_ ;
wire \u_count_l/_19_ ;
wire \u_count_l/_20_ ;
wire \u_count_l/_21_ ;
wire \u_count_l/_22_ ;
wire \u_count_l/_23_ ;
wire \u_count_l/_24_ ;
wire \u_count_l/_25_ ;
wire \u_count_l/_26_ ;
wire \u_count_l/_27_ ;
wire \u_count_l/_28_ ;
wire \u_count_l/_29_ ;
wire \u_count_l/_30_ ;
wire \u_count_l/_31_ ;
wire \u_count_l/_32_ ;
wire \u_count_l/_33_ ;
wire \u_count_l/_34_ ;
wire \u_count_l/_35_ ;
wire \u_count_l/_36_ ;
wire \u_count_l/_37_ ;
wire \u_count_l/_38_ ;
wire \u_count_l/_39_ ;
wire \u_count_l/_40_ ;
wire \u_count_l/_41_ ;
wire \u_count_l/_42_ ;
wire \u_ps2_keyboard/_0000_ ;
wire \u_ps2_keyboard/_0001_ ;
wire \u_ps2_keyboard/_0002_ ;
wire \u_ps2_keyboard/_0003_ ;
wire \u_ps2_keyboard/_0004_ ;
wire \u_ps2_keyboard/_0005_ ;
wire \u_ps2_keyboard/_0006_ ;
wire \u_ps2_keyboard/_0007_ ;
wire \u_ps2_keyboard/_0008_ ;
wire \u_ps2_keyboard/_0009_ ;
wire \u_ps2_keyboard/_0010_ ;
wire \u_ps2_keyboard/_0011_ ;
wire \u_ps2_keyboard/_0012_ ;
wire \u_ps2_keyboard/_0013_ ;
wire \u_ps2_keyboard/_0014_ ;
wire \u_ps2_keyboard/_0015_ ;
wire \u_ps2_keyboard/_0016_ ;
wire \u_ps2_keyboard/_0017_ ;
wire \u_ps2_keyboard/_0018_ ;
wire \u_ps2_keyboard/_0019_ ;
wire \u_ps2_keyboard/_0020_ ;
wire \u_ps2_keyboard/_0021_ ;
wire \u_ps2_keyboard/_0022_ ;
wire \u_ps2_keyboard/_0023_ ;
wire \u_ps2_keyboard/_0024_ ;
wire \u_ps2_keyboard/_0025_ ;
wire \u_ps2_keyboard/_0026_ ;
wire \u_ps2_keyboard/_0027_ ;
wire \u_ps2_keyboard/_0028_ ;
wire \u_ps2_keyboard/_0029_ ;
wire \u_ps2_keyboard/_0030_ ;
wire \u_ps2_keyboard/_0031_ ;
wire \u_ps2_keyboard/_0032_ ;
wire \u_ps2_keyboard/_0033_ ;
wire \u_ps2_keyboard/_0034_ ;
wire \u_ps2_keyboard/_0035_ ;
wire \u_ps2_keyboard/_0036_ ;
wire \u_ps2_keyboard/_0037_ ;
wire \u_ps2_keyboard/_0038_ ;
wire \u_ps2_keyboard/_0039_ ;
wire \u_ps2_keyboard/_0040_ ;
wire \u_ps2_keyboard/_0041_ ;
wire \u_ps2_keyboard/_0042_ ;
wire \u_ps2_keyboard/_0043_ ;
wire \u_ps2_keyboard/_0044_ ;
wire \u_ps2_keyboard/_0045_ ;
wire \u_ps2_keyboard/_0046_ ;
wire \u_ps2_keyboard/_0047_ ;
wire \u_ps2_keyboard/_0048_ ;
wire \u_ps2_keyboard/_0049_ ;
wire \u_ps2_keyboard/_0050_ ;
wire \u_ps2_keyboard/_0051_ ;
wire \u_ps2_keyboard/_0052_ ;
wire \u_ps2_keyboard/_0053_ ;
wire \u_ps2_keyboard/_0054_ ;
wire \u_ps2_keyboard/_0055_ ;
wire \u_ps2_keyboard/_0056_ ;
wire \u_ps2_keyboard/_0057_ ;
wire \u_ps2_keyboard/_0058_ ;
wire \u_ps2_keyboard/_0059_ ;
wire \u_ps2_keyboard/_0060_ ;
wire \u_ps2_keyboard/_0061_ ;
wire \u_ps2_keyboard/_0062_ ;
wire \u_ps2_keyboard/_0063_ ;
wire \u_ps2_keyboard/_0064_ ;
wire \u_ps2_keyboard/_0065_ ;
wire \u_ps2_keyboard/_0066_ ;
wire \u_ps2_keyboard/_0067_ ;
wire \u_ps2_keyboard/_0068_ ;
wire \u_ps2_keyboard/_0069_ ;
wire \u_ps2_keyboard/_0070_ ;
wire \u_ps2_keyboard/_0071_ ;
wire \u_ps2_keyboard/_0072_ ;
wire \u_ps2_keyboard/_0073_ ;
wire \u_ps2_keyboard/_0074_ ;
wire \u_ps2_keyboard/_0075_ ;
wire \u_ps2_keyboard/_0076_ ;
wire \u_ps2_keyboard/_0077_ ;
wire \u_ps2_keyboard/_0078_ ;
wire \u_ps2_keyboard/_0079_ ;
wire \u_ps2_keyboard/_0080_ ;
wire \u_ps2_keyboard/_0081_ ;
wire \u_ps2_keyboard/_0082_ ;
wire \u_ps2_keyboard/_0083_ ;
wire \u_ps2_keyboard/_0084_ ;
wire \u_ps2_keyboard/_0085_ ;
wire \u_ps2_keyboard/_0086_ ;
wire \u_ps2_keyboard/_0087_ ;
wire \u_ps2_keyboard/_0088_ ;
wire \u_ps2_keyboard/_0089_ ;
wire \u_ps2_keyboard/_0090_ ;
wire \u_ps2_keyboard/_0091_ ;
wire \u_ps2_keyboard/_0092_ ;
wire \u_ps2_keyboard/_0093_ ;
wire \u_ps2_keyboard/_0094_ ;
wire \u_ps2_keyboard/_0095_ ;
wire \u_ps2_keyboard/_0096_ ;
wire \u_ps2_keyboard/_0097_ ;
wire \u_ps2_keyboard/_0098_ ;
wire \u_ps2_keyboard/_0099_ ;
wire \u_ps2_keyboard/_0100_ ;
wire \u_ps2_keyboard/_0101_ ;
wire \u_ps2_keyboard/_0102_ ;
wire \u_ps2_keyboard/_0103_ ;
wire \u_ps2_keyboard/_0104_ ;
wire \u_ps2_keyboard/_0105_ ;
wire \u_ps2_keyboard/_0106_ ;
wire \u_ps2_keyboard/_0107_ ;
wire \u_ps2_keyboard/_0108_ ;
wire \u_ps2_keyboard/_0109_ ;
wire \u_ps2_keyboard/_0110_ ;
wire \u_ps2_keyboard/_0111_ ;
wire \u_ps2_keyboard/_0112_ ;
wire \u_ps2_keyboard/_0113_ ;
wire \u_ps2_keyboard/_0114_ ;
wire \u_ps2_keyboard/_0115_ ;
wire \u_ps2_keyboard/_0116_ ;
wire \u_ps2_keyboard/_0117_ ;
wire \u_ps2_keyboard/_0118_ ;
wire \u_ps2_keyboard/_0119_ ;
wire \u_ps2_keyboard/_0120_ ;
wire \u_ps2_keyboard/_0121_ ;
wire \u_ps2_keyboard/_0122_ ;
wire \u_ps2_keyboard/_0123_ ;
wire \u_ps2_keyboard/_0124_ ;
wire \u_ps2_keyboard/_0125_ ;
wire \u_ps2_keyboard/_0126_ ;
wire \u_ps2_keyboard/_0127_ ;
wire \u_ps2_keyboard/_0128_ ;
wire \u_ps2_keyboard/_0129_ ;
wire \u_ps2_keyboard/_0130_ ;
wire \u_ps2_keyboard/_0131_ ;
wire \u_ps2_keyboard/_0132_ ;
wire \u_ps2_keyboard/_0133_ ;
wire \u_ps2_keyboard/_0134_ ;
wire \u_ps2_keyboard/_0135_ ;
wire \u_ps2_keyboard/_0136_ ;
wire \u_ps2_keyboard/_0137_ ;
wire \u_ps2_keyboard/_0138_ ;
wire \u_ps2_keyboard/_0139_ ;
wire \u_ps2_keyboard/_0140_ ;
wire \u_ps2_keyboard/_0141_ ;
wire \u_ps2_keyboard/_0142_ ;
wire \u_ps2_keyboard/_0143_ ;
wire \u_ps2_keyboard/_0144_ ;
wire \u_ps2_keyboard/_0145_ ;
wire \u_ps2_keyboard/_0146_ ;
wire \u_ps2_keyboard/_0147_ ;
wire \u_ps2_keyboard/_0148_ ;
wire \u_ps2_keyboard/_0149_ ;
wire \u_ps2_keyboard/_0150_ ;
wire \u_ps2_keyboard/_0151_ ;
wire \u_ps2_keyboard/_0152_ ;
wire \u_ps2_keyboard/_0153_ ;
wire \u_ps2_keyboard/_0154_ ;
wire \u_ps2_keyboard/_0155_ ;
wire \u_ps2_keyboard/_0156_ ;
wire \u_ps2_keyboard/_0157_ ;
wire \u_ps2_keyboard/_0158_ ;
wire \u_ps2_keyboard/_0159_ ;
wire \u_ps2_keyboard/_0160_ ;
wire \u_ps2_keyboard/_0161_ ;
wire \u_ps2_keyboard/_0162_ ;
wire \u_ps2_keyboard/_0163_ ;
wire \u_ps2_keyboard/_0164_ ;
wire \u_ps2_keyboard/_0165_ ;
wire \u_ps2_keyboard/_0166_ ;
wire \u_ps2_keyboard/_0167_ ;
wire \u_ps2_keyboard/_0168_ ;
wire \u_ps2_keyboard/_0169_ ;
wire \u_ps2_keyboard/_0170_ ;
wire \u_ps2_keyboard/_0171_ ;
wire \u_ps2_keyboard/_0172_ ;
wire \u_ps2_keyboard/_0173_ ;
wire \u_ps2_keyboard/_0174_ ;
wire \u_ps2_keyboard/_0175_ ;
wire \u_ps2_keyboard/_0176_ ;
wire \u_ps2_keyboard/_0177_ ;
wire \u_ps2_keyboard/_0178_ ;
wire \u_ps2_keyboard/_0179_ ;
wire \u_ps2_keyboard/_0180_ ;
wire \u_ps2_keyboard/_0181_ ;
wire \u_ps2_keyboard/_0182_ ;
wire \u_ps2_keyboard/_0183_ ;
wire \u_ps2_keyboard/_0184_ ;
wire \u_ps2_keyboard/_0185_ ;
wire \u_ps2_keyboard/_0186_ ;
wire \u_ps2_keyboard/_0187_ ;
wire \u_ps2_keyboard/_0188_ ;
wire \u_ps2_keyboard/_0189_ ;
wire \u_ps2_keyboard/_0190_ ;
wire \u_ps2_keyboard/_0191_ ;
wire \u_ps2_keyboard/_0192_ ;
wire \u_ps2_keyboard/_0193_ ;
wire \u_ps2_keyboard/_0194_ ;
wire \u_ps2_keyboard/_0195_ ;
wire \u_ps2_keyboard/_0196_ ;
wire \u_ps2_keyboard/_0197_ ;
wire \u_ps2_keyboard/_0198_ ;
wire \u_ps2_keyboard/_0199_ ;
wire \u_ps2_keyboard/_0200_ ;
wire \u_ps2_keyboard/_0201_ ;
wire \u_ps2_keyboard/_0202_ ;
wire \u_ps2_keyboard/_0203_ ;
wire \u_ps2_keyboard/_0204_ ;
wire \u_ps2_keyboard/_0205_ ;
wire \u_ps2_keyboard/_0206_ ;
wire \u_ps2_keyboard/_0207_ ;
wire \u_ps2_keyboard/_0208_ ;
wire \u_ps2_keyboard/_0209_ ;
wire \u_ps2_keyboard/_0210_ ;
wire \u_ps2_keyboard/_0211_ ;
wire \u_ps2_keyboard/_0212_ ;
wire \u_ps2_keyboard/_0213_ ;
wire \u_ps2_keyboard/_0214_ ;
wire \u_ps2_keyboard/_0215_ ;
wire \u_ps2_keyboard/_0216_ ;
wire \u_ps2_keyboard/_0217_ ;
wire \u_ps2_keyboard/_0218_ ;
wire \u_ps2_keyboard/_0219_ ;
wire \u_ps2_keyboard/_0220_ ;
wire \u_ps2_keyboard/_0221_ ;
wire \u_ps2_keyboard/_0222_ ;
wire \u_ps2_keyboard/_0223_ ;
wire \u_ps2_keyboard/_0224_ ;
wire \u_ps2_keyboard/_0225_ ;
wire \u_ps2_keyboard/_0226_ ;
wire \u_ps2_keyboard/_0227_ ;
wire \u_ps2_keyboard/_0228_ ;
wire \u_ps2_keyboard/_0229_ ;
wire \u_ps2_keyboard/_0230_ ;
wire \u_ps2_keyboard/_0231_ ;
wire \u_ps2_keyboard/_0232_ ;
wire \u_ps2_keyboard/_0233_ ;
wire \u_ps2_keyboard/_0234_ ;
wire \u_ps2_keyboard/_0235_ ;
wire \u_ps2_keyboard/_0236_ ;
wire \u_ps2_keyboard/_0237_ ;
wire \u_ps2_keyboard/_0238_ ;
wire \u_ps2_keyboard/_0239_ ;
wire \u_ps2_keyboard/_0240_ ;
wire \u_ps2_keyboard/_0241_ ;
wire \u_ps2_keyboard/_0242_ ;
wire \u_ps2_keyboard/_0243_ ;
wire \u_ps2_keyboard/_0244_ ;
wire \u_ps2_keyboard/_0245_ ;
wire \u_ps2_keyboard/_0246_ ;
wire \u_ps2_keyboard/_0247_ ;
wire \u_ps2_keyboard/_0248_ ;
wire \u_ps2_keyboard/_0249_ ;
wire \u_ps2_keyboard/_0250_ ;
wire \u_ps2_keyboard/_0251_ ;
wire \u_ps2_keyboard/_0252_ ;
wire \u_ps2_keyboard/_0253_ ;
wire \u_ps2_keyboard/_0254_ ;
wire \u_ps2_keyboard/_0255_ ;
wire \u_ps2_keyboard/_0256_ ;
wire \u_ps2_keyboard/_0257_ ;
wire \u_ps2_keyboard/_0258_ ;
wire \u_ps2_keyboard/_0259_ ;
wire \u_ps2_keyboard/_0260_ ;
wire \u_ps2_keyboard/_0261_ ;
wire \u_ps2_keyboard/_0262_ ;
wire \u_ps2_keyboard/_0263_ ;
wire \u_ps2_keyboard/_0264_ ;
wire \u_ps2_keyboard/_0265_ ;
wire \u_ps2_keyboard/_0266_ ;
wire \u_ps2_keyboard/_0267_ ;
wire \u_ps2_keyboard/_0268_ ;
wire \u_ps2_keyboard/_0269_ ;
wire \u_ps2_keyboard/_0270_ ;
wire \u_ps2_keyboard/_0271_ ;
wire \u_ps2_keyboard/_0272_ ;
wire \u_ps2_keyboard/_0273_ ;
wire \u_ps2_keyboard/_0274_ ;
wire \u_ps2_keyboard/_0275_ ;
wire \u_ps2_keyboard/_0276_ ;
wire \u_ps2_keyboard/_0277_ ;
wire \u_ps2_keyboard/_0278_ ;
wire \u_ps2_keyboard/_0279_ ;
wire \u_ps2_keyboard/_0280_ ;
wire \u_ps2_keyboard/_0281_ ;
wire \u_ps2_keyboard/_0282_ ;
wire \u_ps2_keyboard/_0283_ ;
wire \u_ps2_keyboard/_0284_ ;
wire \u_ps2_keyboard/_0285_ ;
wire \u_ps2_keyboard/_0286_ ;
wire \u_ps2_keyboard/_0287_ ;
wire \u_ps2_keyboard/_0288_ ;
wire \u_ps2_keyboard/_0289_ ;
wire \u_ps2_keyboard/_0290_ ;
wire \u_ps2_keyboard/_0291_ ;
wire \u_ps2_keyboard/_0292_ ;
wire \u_ps2_keyboard/_0293_ ;
wire \u_ps2_keyboard/_0294_ ;
wire \u_ps2_keyboard/_0295_ ;
wire \u_ps2_keyboard/_0296_ ;
wire \u_ps2_keyboard/_0297_ ;
wire \u_ps2_keyboard/_0298_ ;
wire \u_ps2_keyboard/_0299_ ;
wire \u_ps2_keyboard/_0300_ ;
wire \u_ps2_keyboard/_0301_ ;
wire \u_ps2_keyboard/_0302_ ;
wire \u_ps2_keyboard/_0303_ ;
wire \u_ps2_keyboard/_0304_ ;
wire \u_ps2_keyboard/_0305_ ;
wire \u_ps2_keyboard/_0306_ ;
wire \u_ps2_keyboard/_0307_ ;
wire \u_ps2_keyboard/_0308_ ;
wire \u_ps2_keyboard/_0309_ ;
wire \u_ps2_keyboard/_0310_ ;
wire \u_ps2_keyboard/_0311_ ;
wire \u_ps2_keyboard/_0312_ ;
wire \u_ps2_keyboard/_0313_ ;
wire \u_ps2_keyboard/_0314_ ;
wire \u_ps2_keyboard/_0315_ ;
wire \u_ps2_keyboard/_0316_ ;
wire \u_ps2_keyboard/_0317_ ;
wire \u_ps2_keyboard/_0318_ ;
wire \u_ps2_keyboard/_0319_ ;
wire \u_ps2_keyboard/_0320_ ;
wire \u_ps2_keyboard/_0321_ ;
wire \u_ps2_keyboard/_0322_ ;
wire \u_ps2_keyboard/_0323_ ;
wire \u_ps2_keyboard/_0324_ ;
wire \u_ps2_keyboard/_0325_ ;
wire \u_ps2_keyboard/_0326_ ;
wire \u_ps2_keyboard/_0327_ ;
wire \u_ps2_keyboard/_0328_ ;
wire \u_ps2_keyboard/_0329_ ;
wire \u_ps2_keyboard/_0330_ ;
wire \u_ps2_keyboard/_0331_ ;
wire \u_ps2_keyboard/_0332_ ;
wire \u_ps2_keyboard/_0333_ ;
wire \u_ps2_keyboard/_0334_ ;
wire \u_ps2_keyboard/_0335_ ;
wire \u_ps2_keyboard/_0336_ ;
wire \u_ps2_keyboard/_0337_ ;
wire \u_ps2_keyboard/_0338_ ;
wire \u_ps2_keyboard/_0339_ ;
wire \u_ps2_keyboard/_0340_ ;
wire \u_ps2_keyboard/_0341_ ;
wire \u_ps2_keyboard/_0342_ ;
wire \u_ps2_keyboard/_0343_ ;
wire \u_ps2_keyboard/_0344_ ;
wire \u_ps2_keyboard/_0345_ ;
wire \u_ps2_keyboard/_0346_ ;
wire \u_ps2_keyboard/_0347_ ;
wire \u_ps2_keyboard/_0348_ ;
wire \u_ps2_keyboard/_0349_ ;
wire \u_ps2_keyboard/_0350_ ;
wire \u_ps2_keyboard/_0351_ ;
wire \u_ps2_keyboard/_0352_ ;
wire \u_ps2_keyboard/_0353_ ;
wire \u_ps2_keyboard/_0354_ ;
wire \u_ps2_keyboard/_0355_ ;
wire \u_ps2_keyboard/_0356_ ;
wire \u_ps2_keyboard/_0357_ ;
wire \u_ps2_keyboard/_0358_ ;
wire \u_ps2_keyboard/_0359_ ;
wire \u_ps2_keyboard/_0360_ ;
wire \u_ps2_keyboard/_0361_ ;
wire \u_ps2_keyboard/_0362_ ;
wire \u_ps2_keyboard/_0363_ ;
wire \u_ps2_keyboard/_0364_ ;
wire \u_ps2_keyboard/_0365_ ;
wire \u_ps2_keyboard/_0366_ ;
wire \u_ps2_keyboard/_0367_ ;
wire \u_ps2_keyboard/_0368_ ;
wire \u_ps2_keyboard/_0369_ ;
wire \u_ps2_keyboard/_0370_ ;
wire \u_ps2_keyboard/_0371_ ;
wire \u_ps2_keyboard/_0372_ ;
wire \u_ps2_keyboard/_0373_ ;
wire \u_ps2_keyboard/_0374_ ;
wire \u_ps2_keyboard/_0375_ ;
wire \u_ps2_keyboard/_0376_ ;
wire \u_ps2_keyboard/_0377_ ;
wire \u_ps2_keyboard/_0378_ ;
wire \u_ps2_keyboard/_0379_ ;
wire \u_ps2_keyboard/_0380_ ;
wire \u_ps2_keyboard/_0381_ ;
wire \u_ps2_keyboard/_0382_ ;
wire \u_ps2_keyboard/_0383_ ;
wire \u_ps2_keyboard/_0384_ ;
wire \u_ps2_keyboard/_0385_ ;
wire \u_ps2_keyboard/_0386_ ;
wire \u_ps2_keyboard/_0387_ ;
wire \u_ps2_keyboard/_0388_ ;
wire \u_ps2_keyboard/_0389_ ;
wire \u_ps2_keyboard/_0390_ ;
wire \u_ps2_keyboard/_0391_ ;
wire \u_ps2_keyboard/_0392_ ;
wire \u_ps2_keyboard/_0393_ ;
wire \u_ps2_keyboard/_0394_ ;
wire \u_ps2_keyboard/_0395_ ;
wire \u_ps2_keyboard/_0396_ ;
wire \u_ps2_keyboard/_0397_ ;
wire \u_ps2_keyboard/_0398_ ;
wire \u_ps2_keyboard/_0399_ ;
wire \u_ps2_keyboard/_0400_ ;
wire \u_ps2_keyboard/_0401_ ;
wire \u_ps2_keyboard/_0402_ ;
wire \u_ps2_keyboard/_0403_ ;
wire \u_ps2_keyboard/_0404_ ;
wire \u_ps2_keyboard/_0405_ ;
wire \u_ps2_keyboard/_0406_ ;
wire \u_ps2_keyboard/_0407_ ;
wire \u_ps2_keyboard/_0408_ ;
wire \u_ps2_keyboard/_0409_ ;
wire \u_ps2_keyboard/_0410_ ;
wire \u_ps2_keyboard/_0411_ ;
wire \u_ps2_keyboard/_0412_ ;
wire \u_ps2_keyboard/_0413_ ;
wire \u_ps2_keyboard/_0414_ ;
wire \u_ps2_keyboard/_0415_ ;
wire \u_ps2_keyboard/_0416_ ;
wire \u_ps2_keyboard/_0417_ ;
wire \u_ps2_keyboard/_0418_ ;
wire \u_ps2_keyboard/_0419_ ;
wire \u_ps2_keyboard/_0420_ ;
wire \u_ps2_keyboard/_0421_ ;
wire \u_ps2_keyboard/_0422_ ;
wire \u_ps2_keyboard/_0423_ ;
wire \u_ps2_keyboard/_0424_ ;
wire \u_ps2_keyboard/_0425_ ;
wire \u_ps2_keyboard/_0426_ ;
wire \u_ps2_keyboard/_0427_ ;
wire \u_ps2_keyboard/_0428_ ;
wire \u_ps2_keyboard/_0429_ ;
wire \u_ps2_keyboard/_0430_ ;
wire \u_ps2_keyboard/_0431_ ;
wire \u_ps2_keyboard/_0432_ ;
wire \u_ps2_keyboard/_0433_ ;
wire \u_ps2_keyboard/_0434_ ;
wire \u_ps2_keyboard/_0435_ ;
wire \u_ps2_keyboard/_0436_ ;
wire \u_ps2_keyboard/_0437_ ;
wire \u_ps2_keyboard/_0438_ ;
wire \u_ps2_keyboard/_0439_ ;
wire \u_ps2_keyboard/_0440_ ;
wire \u_ps2_keyboard/_0441_ ;
wire \u_ps2_keyboard/_0442_ ;
wire \u_ps2_keyboard/_0443_ ;
wire \u_ps2_keyboard/_0444_ ;
wire \u_ps2_keyboard/_0445_ ;
wire \u_ps2_keyboard/_0446_ ;
wire \u_ps2_keyboard/_0447_ ;
wire \u_ps2_keyboard/_0448_ ;
wire \u_ps2_keyboard/_0449_ ;
wire \u_ps2_keyboard/_0450_ ;
wire \u_ps2_keyboard/_0451_ ;
wire \u_ps2_keyboard/_0452_ ;
wire \u_ps2_keyboard/_0453_ ;
wire \u_ps2_keyboard/_0454_ ;
wire \u_ps2_keyboard/_0455_ ;
wire \u_ps2_keyboard/_0456_ ;
wire \u_ps2_keyboard/_0457_ ;
wire \u_ps2_keyboard/_0458_ ;
wire \u_ps2_keyboard/_0459_ ;
wire \u_ps2_keyboard/_0460_ ;
wire \u_ps2_keyboard/_0461_ ;
wire \u_ps2_keyboard/_0462_ ;
wire \u_ps2_keyboard/_0463_ ;
wire \u_ps2_keyboard/_0464_ ;
wire \u_ps2_keyboard/_0465_ ;
wire \u_ps2_keyboard/_0466_ ;
wire \u_ps2_keyboard/_0467_ ;
wire \u_ps2_keyboard/_0468_ ;
wire \u_ps2_keyboard/_0469_ ;
wire \u_ps2_keyboard/_0470_ ;
wire \u_ps2_keyboard/_0471_ ;
wire \u_ps2_keyboard/_0472_ ;
wire \u_ps2_keyboard/_0473_ ;
wire \u_ps2_keyboard/_0474_ ;
wire \u_ps2_keyboard/_0475_ ;
wire \u_ps2_keyboard/_0476_ ;
wire \u_ps2_keyboard/_0477_ ;
wire \u_ps2_keyboard/_0478_ ;
wire \u_ps2_keyboard/_0479_ ;
wire \u_ps2_keyboard/_0480_ ;
wire \u_ps2_keyboard/_0481_ ;
wire \u_ps2_keyboard/_0482_ ;
wire \u_ps2_keyboard/_0483_ ;
wire \u_ps2_keyboard/_0484_ ;
wire \u_ps2_keyboard/_0485_ ;
wire \u_ps2_keyboard/_0486_ ;
wire \u_ps2_keyboard/_0487_ ;
wire \u_ps2_keyboard/_0488_ ;
wire \u_ps2_keyboard/_0489_ ;
wire \u_ps2_keyboard/_0490_ ;
wire \u_ps2_keyboard/_0491_ ;
wire \u_ps2_keyboard/_0492_ ;
wire \u_ps2_keyboard/_0493_ ;
wire \u_ps2_keyboard/_0494_ ;
wire \u_ps2_keyboard/_0495_ ;
wire \u_ps2_keyboard/_0496_ ;
wire \u_ps2_keyboard/_0497_ ;
wire \u_ps2_keyboard/_0498_ ;
wire \u_ps2_keyboard/_0499_ ;
wire \u_ps2_keyboard/_0500_ ;
wire \u_ps2_keyboard/_0501_ ;
wire \u_ps2_keyboard/_0502_ ;
wire \u_ps2_keyboard/_0503_ ;
wire \u_ps2_keyboard/_0504_ ;
wire \u_ps2_keyboard/_0505_ ;
wire \u_ps2_keyboard/_0506_ ;
wire \u_ps2_keyboard/_0507_ ;
wire \u_ps2_keyboard/_0508_ ;
wire \u_ps2_keyboard/_0509_ ;
wire \u_ps2_keyboard/_0510_ ;
wire \u_ps2_keyboard/_0511_ ;
wire \u_ps2_keyboard/_0512_ ;
wire \u_ps2_keyboard/_0513_ ;
wire \u_ps2_keyboard/_0514_ ;
wire \u_ps2_keyboard/_0515_ ;
wire \u_ps2_keyboard/_0516_ ;
wire \u_ps2_keyboard/_0517_ ;
wire \u_ps2_keyboard/_0518_ ;
wire \u_ps2_keyboard/_0519_ ;
wire \u_ps2_keyboard/_0520_ ;
wire \u_ps2_keyboard/_0521_ ;
wire \u_ps2_keyboard/_0522_ ;
wire \u_ps2_keyboard/_0523_ ;
wire \u_ps2_keyboard/_0524_ ;
wire \u_ps2_keyboard/_0525_ ;
wire \u_ps2_keyboard/_0526_ ;
wire \u_ps2_keyboard/_0527_ ;
wire \u_ps2_keyboard/fifo[0][0] ;
wire \u_ps2_keyboard/fifo[0][1] ;
wire \u_ps2_keyboard/fifo[0][2] ;
wire \u_ps2_keyboard/fifo[0][3] ;
wire \u_ps2_keyboard/fifo[0][4] ;
wire \u_ps2_keyboard/fifo[0][5] ;
wire \u_ps2_keyboard/fifo[0][6] ;
wire \u_ps2_keyboard/fifo[0][7] ;
wire \u_ps2_keyboard/fifo[1][0] ;
wire \u_ps2_keyboard/fifo[1][1] ;
wire \u_ps2_keyboard/fifo[1][2] ;
wire \u_ps2_keyboard/fifo[1][3] ;
wire \u_ps2_keyboard/fifo[1][4] ;
wire \u_ps2_keyboard/fifo[1][5] ;
wire \u_ps2_keyboard/fifo[1][6] ;
wire \u_ps2_keyboard/fifo[1][7] ;
wire \u_ps2_keyboard/fifo[2][0] ;
wire \u_ps2_keyboard/fifo[2][1] ;
wire \u_ps2_keyboard/fifo[2][2] ;
wire \u_ps2_keyboard/fifo[2][3] ;
wire \u_ps2_keyboard/fifo[2][4] ;
wire \u_ps2_keyboard/fifo[2][5] ;
wire \u_ps2_keyboard/fifo[2][6] ;
wire \u_ps2_keyboard/fifo[2][7] ;
wire \u_ps2_keyboard/fifo[3][0] ;
wire \u_ps2_keyboard/fifo[3][1] ;
wire \u_ps2_keyboard/fifo[3][2] ;
wire \u_ps2_keyboard/fifo[3][3] ;
wire \u_ps2_keyboard/fifo[3][4] ;
wire \u_ps2_keyboard/fifo[3][5] ;
wire \u_ps2_keyboard/fifo[3][6] ;
wire \u_ps2_keyboard/fifo[3][7] ;
wire \u_ps2_keyboard/fifo[4][0] ;
wire \u_ps2_keyboard/fifo[4][1] ;
wire \u_ps2_keyboard/fifo[4][2] ;
wire \u_ps2_keyboard/fifo[4][3] ;
wire \u_ps2_keyboard/fifo[4][4] ;
wire \u_ps2_keyboard/fifo[4][5] ;
wire \u_ps2_keyboard/fifo[4][6] ;
wire \u_ps2_keyboard/fifo[4][7] ;
wire \u_ps2_keyboard/fifo[5][0] ;
wire \u_ps2_keyboard/fifo[5][1] ;
wire \u_ps2_keyboard/fifo[5][2] ;
wire \u_ps2_keyboard/fifo[5][3] ;
wire \u_ps2_keyboard/fifo[5][4] ;
wire \u_ps2_keyboard/fifo[5][5] ;
wire \u_ps2_keyboard/fifo[5][6] ;
wire \u_ps2_keyboard/fifo[5][7] ;
wire \u_ps2_keyboard/fifo[6][0] ;
wire \u_ps2_keyboard/fifo[6][1] ;
wire \u_ps2_keyboard/fifo[6][2] ;
wire \u_ps2_keyboard/fifo[6][3] ;
wire \u_ps2_keyboard/fifo[6][4] ;
wire \u_ps2_keyboard/fifo[6][5] ;
wire \u_ps2_keyboard/fifo[6][6] ;
wire \u_ps2_keyboard/fifo[6][7] ;
wire \u_ps2_keyboard/fifo[7][0] ;
wire \u_ps2_keyboard/fifo[7][1] ;
wire \u_ps2_keyboard/fifo[7][2] ;
wire \u_ps2_keyboard/fifo[7][3] ;
wire \u_ps2_keyboard/fifo[7][4] ;
wire \u_ps2_keyboard/fifo[7][5] ;
wire \u_ps2_keyboard/fifo[7][6] ;
wire \u_ps2_keyboard/fifo[7][7] ;
wire \u_rom/_000_ ;
wire \u_rom/_001_ ;
wire \u_rom/_002_ ;
wire \u_rom/_003_ ;
wire \u_rom/_004_ ;
wire \u_rom/_005_ ;
wire \u_rom/_006_ ;
wire \u_rom/_007_ ;
wire \u_rom/_008_ ;
wire \u_rom/_009_ ;
wire \u_rom/_010_ ;
wire \u_rom/_011_ ;
wire \u_rom/_012_ ;
wire \u_rom/_013_ ;
wire \u_rom/_014_ ;
wire \u_rom/_015_ ;
wire \u_rom/_016_ ;
wire \u_rom/_017_ ;
wire \u_rom/_018_ ;
wire \u_rom/_019_ ;
wire \u_rom/_020_ ;
wire \u_rom/_021_ ;
wire \u_rom/_022_ ;
wire \u_rom/_023_ ;
wire \u_rom/_024_ ;
wire \u_rom/_025_ ;
wire \u_rom/_026_ ;
wire \u_rom/_027_ ;
wire \u_rom/_028_ ;
wire \u_rom/_029_ ;
wire \u_rom/_030_ ;
wire \u_rom/_031_ ;
wire \u_rom/_032_ ;
wire \u_rom/_033_ ;
wire \u_rom/_034_ ;
wire \u_rom/_035_ ;
wire \u_rom/_036_ ;
wire \u_rom/_037_ ;
wire \u_rom/_038_ ;
wire \u_rom/_039_ ;
wire \u_rom/_040_ ;
wire \u_rom/_041_ ;
wire \u_rom/_042_ ;
wire \u_rom/_043_ ;
wire \u_rom/_044_ ;
wire \u_rom/_045_ ;
wire \u_rom/_046_ ;
wire \u_rom/_047_ ;
wire \u_rom/_048_ ;
wire \u_rom/_049_ ;
wire \u_scan_code_h/_00_ ;
wire \u_scan_code_h/_01_ ;
wire \u_scan_code_h/_02_ ;
wire \u_scan_code_h/_03_ ;
wire \u_scan_code_h/_04_ ;
wire \u_scan_code_h/_05_ ;
wire \u_scan_code_h/_06_ ;
wire \u_scan_code_h/_07_ ;
wire \u_scan_code_h/_08_ ;
wire \u_scan_code_h/_09_ ;
wire \u_scan_code_h/_10_ ;
wire \u_scan_code_h/_11_ ;
wire \u_scan_code_h/_12_ ;
wire \u_scan_code_h/_13_ ;
wire \u_scan_code_h/_14_ ;
wire \u_scan_code_h/_15_ ;
wire \u_scan_code_h/_16_ ;
wire \u_scan_code_h/_17_ ;
wire \u_scan_code_h/_18_ ;
wire \u_scan_code_h/_19_ ;
wire \u_scan_code_h/_20_ ;
wire \u_scan_code_h/_21_ ;
wire \u_scan_code_h/_22_ ;
wire \u_scan_code_h/_23_ ;
wire \u_scan_code_h/_24_ ;
wire \u_scan_code_h/_25_ ;
wire \u_scan_code_h/_26_ ;
wire \u_scan_code_h/_27_ ;
wire \u_scan_code_h/_28_ ;
wire \u_scan_code_h/_29_ ;
wire \u_scan_code_h/_30_ ;
wire \u_scan_code_h/_31_ ;
wire \u_scan_code_h/_32_ ;
wire \u_scan_code_h/_33_ ;
wire \u_scan_code_h/_34_ ;
wire \u_scan_code_h/_35_ ;
wire \u_scan_code_h/_36_ ;
wire \u_scan_code_h/_37_ ;
wire \u_scan_code_h/_38_ ;
wire \u_scan_code_h/_39_ ;
wire \u_scan_code_h/_40_ ;
wire \u_scan_code_h/_41_ ;
wire \u_scan_code_h/_42_ ;
wire \u_scan_code_l/_00_ ;
wire \u_scan_code_l/_01_ ;
wire \u_scan_code_l/_02_ ;
wire \u_scan_code_l/_03_ ;
wire \u_scan_code_l/_04_ ;
wire \u_scan_code_l/_05_ ;
wire \u_scan_code_l/_06_ ;
wire \u_scan_code_l/_07_ ;
wire \u_scan_code_l/_08_ ;
wire \u_scan_code_l/_09_ ;
wire \u_scan_code_l/_10_ ;
wire \u_scan_code_l/_11_ ;
wire \u_scan_code_l/_12_ ;
wire \u_scan_code_l/_13_ ;
wire \u_scan_code_l/_14_ ;
wire \u_scan_code_l/_15_ ;
wire \u_scan_code_l/_16_ ;
wire \u_scan_code_l/_17_ ;
wire \u_scan_code_l/_18_ ;
wire \u_scan_code_l/_19_ ;
wire \u_scan_code_l/_20_ ;
wire \u_scan_code_l/_21_ ;
wire \u_scan_code_l/_22_ ;
wire \u_scan_code_l/_23_ ;
wire \u_scan_code_l/_24_ ;
wire \u_scan_code_l/_25_ ;
wire \u_scan_code_l/_26_ ;
wire \u_scan_code_l/_27_ ;
wire \u_scan_code_l/_28_ ;
wire \u_scan_code_l/_29_ ;
wire \u_scan_code_l/_30_ ;
wire \u_scan_code_l/_31_ ;
wire \u_scan_code_l/_32_ ;
wire \u_scan_code_l/_33_ ;
wire \u_scan_code_l/_34_ ;
wire \u_scan_code_l/_35_ ;
wire \u_scan_code_l/_36_ ;
wire \u_scan_code_l/_37_ ;
wire \u_scan_code_l/_38_ ;
wire \u_scan_code_l/_39_ ;
wire \u_scan_code_l/_40_ ;
wire \u_scan_code_l/_41_ ;
wire \u_scan_code_l/_42_ ;
wire rst_n ;
wire clk ;
wire ps2_data ;
wire overflow ;
wire ps2_clk ;
wire [7:0] ascii_code ;
wire [7:0] count ;
wire [7:0] scan_code ;
wire [7:0] scan_code_buf ;
wire [2:0] state ;
wire [9:0] \u_ps2_keyboard/buffer ;
wire [3:0] \u_ps2_keyboard/count ;
wire [2:0] \u_ps2_keyboard/ps2_clk_sync ;
wire [2:0] \u_ps2_keyboard/r_ptr ;
wire [2:0] \u_ps2_keyboard/w_ptr ;
wire [15:0] ascii_seg ;
wire [15:0] count_seg ;
wire [15:0] scan_code_seg ;


AND2_X4 _143_ ( .A1(_120_ ), .A2(_119_ ), .ZN(_085_ ) );
AND3_X2 _144_ ( .A1(_085_ ), .A2(_122_ ), .A3(_121_ ), .ZN(_086_ ) );
NOR4_X4 _145_ ( .A1(_116_ ), .A2(_115_ ), .A3(_118_ ), .A4(_117_ ), .ZN(_087_ ) );
NAND4_X1 _146_ ( .A1(_086_ ), .A2(_114_ ), .A3(_087_ ), .A4(_113_ ), .ZN(_088_ ) );
NAND2_X1 _147_ ( .A1(_114_ ), .A2(_113_ ), .ZN(_089_ ) );
OAI22_X1 _148_ ( .A1(_088_ ), .A2(_053_ ), .B1(_052_ ), .B2(_089_ ), .ZN(_046_ ) );
AND2_X2 _149_ ( .A1(_086_ ), .A2(_087_ ), .ZN(_090_ ) );
AND2_X2 _150_ ( .A1(_090_ ), .A2(_113_ ), .ZN(_091_ ) );
INV_X1 _151_ ( .A(_114_ ), .ZN(_092_ ) );
OR3_X2 _152_ ( .A1(_091_ ), .A2(_092_ ), .A3(_053_ ), .ZN(_093_ ) );
OAI21_X1 _153_ ( .A(_093_ ), .B1(_054_ ), .B2(_089_ ), .ZN(_047_ ) );
NOR3_X1 _154_ ( .A1(_092_ ), .A2(_131_ ), .A3(_065_ ), .ZN(_094_ ) );
AOI21_X1 _155_ ( .A(_094_ ), .B1(_114_ ), .B2(_113_ ), .ZN(_045_ ) );
AOI21_X1 _156_ ( .A(_053_ ), .B1(_086_ ), .B2(_087_ ), .ZN(_066_ ) );
MUX2_X1 _157_ ( .A(_123_ ), .B(_115_ ), .S(_113_ ), .Z(_095_ ) );
AND2_X1 _158_ ( .A1(_095_ ), .A2(_114_ ), .ZN(_037_ ) );
MUX2_X1 _159_ ( .A(_124_ ), .B(_116_ ), .S(_113_ ), .Z(_096_ ) );
AND2_X1 _160_ ( .A1(_096_ ), .A2(_114_ ), .ZN(_038_ ) );
MUX2_X1 _161_ ( .A(_125_ ), .B(_117_ ), .S(_113_ ), .Z(_097_ ) );
AND2_X1 _162_ ( .A1(_097_ ), .A2(_114_ ), .ZN(_039_ ) );
MUX2_X1 _163_ ( .A(_126_ ), .B(_118_ ), .S(_113_ ), .Z(_098_ ) );
AND2_X1 _164_ ( .A1(_098_ ), .A2(_114_ ), .ZN(_040_ ) );
MUX2_X1 _165_ ( .A(_127_ ), .B(_119_ ), .S(_113_ ), .Z(_099_ ) );
AND2_X1 _166_ ( .A1(_099_ ), .A2(_114_ ), .ZN(_041_ ) );
MUX2_X1 _167_ ( .A(_128_ ), .B(_120_ ), .S(_113_ ), .Z(_100_ ) );
AND2_X1 _168_ ( .A1(_100_ ), .A2(_114_ ), .ZN(_042_ ) );
MUX2_X1 _169_ ( .A(_129_ ), .B(_121_ ), .S(_113_ ), .Z(_101_ ) );
AND2_X1 _170_ ( .A1(_101_ ), .A2(_114_ ), .ZN(_043_ ) );
MUX2_X1 _171_ ( .A(_130_ ), .B(_122_ ), .S(_113_ ), .Z(_102_ ) );
AND2_X1 _172_ ( .A1(_102_ ), .A2(_114_ ), .ZN(_044_ ) );
OAI21_X1 _173_ ( .A(_114_ ), .B1(_065_ ), .B2(_058_ ), .ZN(_103_ ) );
AOI21_X1 _174_ ( .A(_103_ ), .B1(_065_ ), .B2(_058_ ), .ZN(_029_ ) );
INV_X32 _175_ ( .A(_065_ ), .ZN(_104_ ) );
AND2_X4 _176_ ( .A1(_058_ ), .A2(_059_ ), .ZN(_105_ ) );
INV_X4 _177_ ( .A(_105_ ), .ZN(_106_ ) );
OR2_X1 _178_ ( .A1(_058_ ), .A2(_059_ ), .ZN(_107_ ) );
AOI21_X1 _179_ ( .A(_104_ ), .B1(_106_ ), .B2(_107_ ), .ZN(_108_ ) );
AOI211_X4 _180_ ( .A(_092_ ), .B(_108_ ), .C1(_104_ ), .C2(_055_ ), .ZN(_030_ ) );
AND2_X1 _181_ ( .A1(_105_ ), .A2(_060_ ), .ZN(_109_ ) );
AND2_X1 _182_ ( .A1(_109_ ), .A2(_065_ ), .ZN(_110_ ) );
AND2_X1 _183_ ( .A1(_104_ ), .A2(_056_ ), .ZN(_111_ ) );
NOR3_X1 _184_ ( .A1(_105_ ), .A2(_104_ ), .A3(_060_ ), .ZN(_112_ ) );
NOR4_X1 _185_ ( .A1(_110_ ), .A2(_092_ ), .A3(_111_ ), .A4(_112_ ), .ZN(_031_ ) );
XNOR2_X1 _186_ ( .A(_110_ ), .B(_057_ ), .ZN(_067_ ) );
AND2_X1 _187_ ( .A1(_067_ ), .A2(_114_ ), .ZN(_032_ ) );
NAND2_X4 _188_ ( .A1(_060_ ), .A2(_061_ ), .ZN(_068_ ) );
NOR3_X4 _189_ ( .A1(_106_ ), .A2(_104_ ), .A3(_068_ ), .ZN(_069_ ) );
AND2_X1 _190_ ( .A1(_069_ ), .A2(_062_ ), .ZN(_070_ ) );
NOR2_X4 _191_ ( .A1(_106_ ), .A2(_068_ ), .ZN(_071_ ) );
NOR3_X1 _192_ ( .A1(_071_ ), .A2(_104_ ), .A3(_062_ ), .ZN(_072_ ) );
AND2_X1 _193_ ( .A1(_104_ ), .A2(_048_ ), .ZN(_073_ ) );
NOR4_X1 _194_ ( .A1(_070_ ), .A2(_072_ ), .A3(_092_ ), .A4(_073_ ), .ZN(_033_ ) );
OR2_X1 _195_ ( .A1(_070_ ), .A2(_049_ ), .ZN(_074_ ) );
NAND4_X1 _196_ ( .A1(_071_ ), .A2(_065_ ), .A3(_062_ ), .A4(_049_ ), .ZN(_075_ ) );
AOI21_X1 _197_ ( .A(_092_ ), .B1(_074_ ), .B2(_075_ ), .ZN(_034_ ) );
AND2_X1 _198_ ( .A1(_062_ ), .A2(_063_ ), .ZN(_076_ ) );
AND2_X4 _199_ ( .A1(_071_ ), .A2(_076_ ), .ZN(_077_ ) );
OR2_X2 _200_ ( .A1(_077_ ), .A2(_064_ ), .ZN(_078_ ) );
NAND3_X1 _201_ ( .A1(_071_ ), .A2(_064_ ), .A3(_076_ ), .ZN(_079_ ) );
AOI21_X2 _202_ ( .A(_104_ ), .B1(_078_ ), .B2(_079_ ), .ZN(_080_ ) );
AOI211_X2 _203_ ( .A(_092_ ), .B(_080_ ), .C1(_104_ ), .C2(_050_ ), .ZN(_035_ ) );
AND3_X2 _204_ ( .A1(_069_ ), .A2(_064_ ), .A3(_076_ ), .ZN(_081_ ) );
INV_X1 _205_ ( .A(_081_ ), .ZN(_082_ ) );
OR2_X2 _206_ ( .A1(_082_ ), .A2(_051_ ), .ZN(_083_ ) );
AOI21_X1 _207_ ( .A(_092_ ), .B1(_082_ ), .B2(_051_ ), .ZN(_084_ ) );
AND2_X1 _208_ ( .A1(_083_ ), .A2(_084_ ), .ZN(_036_ ) );
LOGIC1_X1 _209_ ( .Z(_141_ ) );
LOGIC0_X1 _210_ ( .Z(_142_ ) );
BUF_X1 _211_ ( .A(count_en ), .Z(\state [1] ) );
BUF_X1 _212_ ( .A(rst_n ), .Z(_114_ ) );
BUF_X1 _213_ ( .A(ready ), .Z(_113_ ) );
BUF_X1 _214_ ( .A(\scan_code [1] ), .Z(_116_ ) );
BUF_X1 _215_ ( .A(\scan_code [0] ), .Z(_115_ ) );
BUF_X1 _216_ ( .A(\scan_code [3] ), .Z(_118_ ) );
BUF_X1 _217_ ( .A(\scan_code [2] ), .Z(_117_ ) );
BUF_X1 _218_ ( .A(\scan_code [5] ), .Z(_120_ ) );
BUF_X1 _219_ ( .A(\scan_code [4] ), .Z(_119_ ) );
BUF_X1 _220_ ( .A(\scan_code [7] ), .Z(_122_ ) );
BUF_X1 _221_ ( .A(\scan_code [6] ), .Z(_121_ ) );
BUF_X1 _222_ ( .A(_024_ ), .Z(_053_ ) );
BUF_X1 _223_ ( .A(_023_ ), .Z(_052_ ) );
BUF_X1 _224_ ( .A(_046_ ), .Z(_017_ ) );
BUF_X1 _225_ ( .A(_025_ ), .Z(_054_ ) );
BUF_X1 _226_ ( .A(_047_ ), .Z(_018_ ) );
BUF_X1 _227_ ( .A(\state [0] ), .Z(_131_ ) );
BUF_X1 _228_ ( .A(count_en ), .Z(_065_ ) );
BUF_X1 _229_ ( .A(_045_ ), .Z(_016_ ) );
BUF_X1 _230_ ( .A(_066_ ), .Z(display_en ) );
BUF_X1 _231_ ( .A(\scan_code_buf [0] ), .Z(_123_ ) );
BUF_X1 _232_ ( .A(_037_ ), .Z(_008_ ) );
BUF_X1 _233_ ( .A(\scan_code_buf [1] ), .Z(_124_ ) );
BUF_X1 _234_ ( .A(_038_ ), .Z(_009_ ) );
BUF_X1 _235_ ( .A(\scan_code_buf [2] ), .Z(_125_ ) );
BUF_X1 _236_ ( .A(_039_ ), .Z(_010_ ) );
BUF_X1 _237_ ( .A(\scan_code_buf [3] ), .Z(_126_ ) );
BUF_X1 _238_ ( .A(_040_ ), .Z(_011_ ) );
BUF_X1 _239_ ( .A(\scan_code_buf [4] ), .Z(_127_ ) );
BUF_X1 _240_ ( .A(_041_ ), .Z(_012_ ) );
BUF_X1 _241_ ( .A(\scan_code_buf [5] ), .Z(_128_ ) );
BUF_X1 _242_ ( .A(_042_ ), .Z(_013_ ) );
BUF_X1 _243_ ( .A(\scan_code_buf [6] ), .Z(_129_ ) );
BUF_X1 _244_ ( .A(_043_ ), .Z(_014_ ) );
BUF_X1 _245_ ( .A(\scan_code_buf [7] ), .Z(_130_ ) );
BUF_X1 _246_ ( .A(_044_ ), .Z(_015_ ) );
BUF_X1 _247_ ( .A(\count [0] ), .Z(_058_ ) );
BUF_X1 _248_ ( .A(_029_ ), .Z(_000_ ) );
BUF_X1 _249_ ( .A(\count [1] ), .Z(_059_ ) );
BUF_X1 _250_ ( .A(_026_ ), .Z(_055_ ) );
BUF_X1 _251_ ( .A(_030_ ), .Z(_001_ ) );
BUF_X1 _252_ ( .A(\count [2] ), .Z(_060_ ) );
BUF_X1 _253_ ( .A(_027_ ), .Z(_056_ ) );
BUF_X1 _254_ ( .A(_031_ ), .Z(_002_ ) );
BUF_X1 _255_ ( .A(_028_ ), .Z(_057_ ) );
BUF_X1 _256_ ( .A(_032_ ), .Z(_003_ ) );
BUF_X1 _257_ ( .A(\count [3] ), .Z(_061_ ) );
BUF_X1 _258_ ( .A(\count [4] ), .Z(_062_ ) );
BUF_X1 _259_ ( .A(_019_ ), .Z(_048_ ) );
BUF_X1 _260_ ( .A(_033_ ), .Z(_004_ ) );
BUF_X1 _261_ ( .A(_020_ ), .Z(_049_ ) );
BUF_X1 _262_ ( .A(_034_ ), .Z(_005_ ) );
BUF_X1 _263_ ( .A(\count [5] ), .Z(_063_ ) );
BUF_X1 _264_ ( .A(\count [6] ), .Z(_064_ ) );
BUF_X1 _265_ ( .A(_021_ ), .Z(_050_ ) );
BUF_X1 _266_ ( .A(_035_ ), .Z(_006_ ) );
BUF_X1 _267_ ( .A(_022_ ), .Z(_051_ ) );
BUF_X1 _268_ ( .A(_036_ ), .Z(_007_ ) );
DFF_X1 _269_ ( .D(_016_ ), .CK(clk ), .Q(\state [0] ), .QN(_025_ ) );
DFF_X1 _270_ ( .D(_017_ ), .CK(clk ), .Q(count_en ), .QN(_023_ ) );
DFF_X1 _271_ ( .D(_018_ ), .CK(clk ), .Q(\state [2] ), .QN(_024_ ) );
DFF_X1 _272_ ( .D(_000_ ), .CK(clk ), .Q(\count [0] ), .QN(_132_ ) );
DFF_X1 _273_ ( .D(_001_ ), .CK(clk ), .Q(\count [1] ), .QN(_026_ ) );
DFF_X1 _274_ ( .D(_002_ ), .CK(clk ), .Q(\count [2] ), .QN(_027_ ) );
DFF_X1 _275_ ( .D(_003_ ), .CK(clk ), .Q(\count [3] ), .QN(_028_ ) );
DFF_X1 _276_ ( .D(_004_ ), .CK(clk ), .Q(\count [4] ), .QN(_019_ ) );
DFF_X1 _277_ ( .D(_005_ ), .CK(clk ), .Q(\count [5] ), .QN(_020_ ) );
DFF_X1 _278_ ( .D(_006_ ), .CK(clk ), .Q(\count [6] ), .QN(_021_ ) );
DFF_X1 _279_ ( .D(_007_ ), .CK(clk ), .Q(\count [7] ), .QN(_022_ ) );
DFF_X1 _280_ ( .D(_008_ ), .CK(clk ), .Q(\scan_code_buf [0] ), .QN(_133_ ) );
DFF_X1 _281_ ( .D(_009_ ), .CK(clk ), .Q(\scan_code_buf [1] ), .QN(_134_ ) );
DFF_X1 _282_ ( .D(_010_ ), .CK(clk ), .Q(\scan_code_buf [2] ), .QN(_135_ ) );
DFF_X1 _283_ ( .D(_011_ ), .CK(clk ), .Q(\scan_code_buf [3] ), .QN(_136_ ) );
DFF_X1 _284_ ( .D(_012_ ), .CK(clk ), .Q(\scan_code_buf [4] ), .QN(_137_ ) );
DFF_X1 _285_ ( .D(_013_ ), .CK(clk ), .Q(\scan_code_buf [5] ), .QN(_138_ ) );
DFF_X1 _286_ ( .D(_014_ ), .CK(clk ), .Q(\scan_code_buf [6] ), .QN(_139_ ) );
DFF_X1 _287_ ( .D(_015_ ), .CK(clk ), .Q(\scan_code_buf [7] ), .QN(_140_ ) );
NOR2_X4 \u_ascii_h/_43_ ( .A1(\u_ascii_h/_01_ ), .A2(\u_ascii_h/_00_ ), .ZN(\u_ascii_h/_05_ ) );
INV_X2 \u_ascii_h/_44_ ( .A(\u_ascii_h/_05_ ), .ZN(\u_ascii_h/_06_ ) );
INV_X4 \u_ascii_h/_45_ ( .A(\u_ascii_h/_02_ ), .ZN(\u_ascii_h/_07_ ) );
NOR2_X2 \u_ascii_h/_46_ ( .A1(\u_ascii_h/_07_ ), .A2(\u_ascii_h/_03_ ), .ZN(\u_ascii_h/_08_ ) );
INV_X16 \u_ascii_h/_47_ ( .A(\u_ascii_h/_03_ ), .ZN(\u_ascii_h/_09_ ) );
NOR2_X2 \u_ascii_h/_48_ ( .A1(\u_ascii_h/_09_ ), .A2(\u_ascii_h/_02_ ), .ZN(\u_ascii_h/_10_ ) );
OR3_X4 \u_ascii_h/_49_ ( .A1(\u_ascii_h/_06_ ), .A2(\u_ascii_h/_08_ ), .A3(\u_ascii_h/_10_ ), .ZN(\u_ascii_h/_11_ ) );
INV_X32 \u_ascii_h/_50_ ( .A(\u_ascii_h/_00_ ), .ZN(\u_ascii_h/_12_ ) );
NOR2_X2 \u_ascii_h/_51_ ( .A1(\u_ascii_h/_12_ ), .A2(\u_ascii_h/_01_ ), .ZN(\u_ascii_h/_13_ ) );
NOR2_X4 \u_ascii_h/_52_ ( .A1(\u_ascii_h/_03_ ), .A2(\u_ascii_h/_02_ ), .ZN(\u_ascii_h/_14_ ) );
AND2_X1 \u_ascii_h/_53_ ( .A1(\u_ascii_h/_13_ ), .A2(\u_ascii_h/_14_ ), .ZN(\u_ascii_h/_15_ ) );
INV_X1 \u_ascii_h/_54_ ( .A(\u_ascii_h/_15_ ), .ZN(\u_ascii_h/_16_ ) );
INV_X1 \u_ascii_h/_55_ ( .A(\u_ascii_h/_04_ ), .ZN(\u_ascii_h/_17_ ) );
AND2_X4 \u_ascii_h/_56_ ( .A1(\u_ascii_h/_01_ ), .A2(\u_ascii_h/_00_ ), .ZN(\u_ascii_h/_18_ ) );
AOI21_X1 \u_ascii_h/_57_ ( .A(\u_ascii_h/_17_ ), .B1(\u_ascii_h/_08_ ), .B2(\u_ascii_h/_18_ ), .ZN(\u_ascii_h/_19_ ) );
NAND3_X1 \u_ascii_h/_58_ ( .A1(\u_ascii_h/_11_ ), .A2(\u_ascii_h/_16_ ), .A3(\u_ascii_h/_19_ ), .ZN(\u_ascii_h/_35_ ) );
NAND2_X1 \u_ascii_h/_59_ ( .A1(\u_ascii_h/_06_ ), .A2(\u_ascii_h/_14_ ), .ZN(\u_ascii_h/_20_ ) );
AND2_X2 \u_ascii_h/_60_ ( .A1(\u_ascii_h/_03_ ), .A2(\u_ascii_h/_02_ ), .ZN(\u_ascii_h/_21_ ) );
NAND2_X1 \u_ascii_h/_61_ ( .A1(\u_ascii_h/_13_ ), .A2(\u_ascii_h/_21_ ), .ZN(\u_ascii_h/_22_ ) );
NAND3_X1 \u_ascii_h/_62_ ( .A1(\u_ascii_h/_19_ ), .A2(\u_ascii_h/_20_ ), .A3(\u_ascii_h/_22_ ), .ZN(\u_ascii_h/_36_ ) );
NOR3_X1 \u_ascii_h/_63_ ( .A1(\u_ascii_h/_07_ ), .A2(\u_ascii_h/_03_ ), .A3(\u_ascii_h/_01_ ), .ZN(\u_ascii_h/_23_ ) );
AOI21_X1 \u_ascii_h/_64_ ( .A(\u_ascii_h/_23_ ), .B1(\u_ascii_h/_08_ ), .B2(\u_ascii_h/_18_ ), .ZN(\u_ascii_h/_24_ ) );
NAND3_X1 \u_ascii_h/_65_ ( .A1(\u_ascii_h/_09_ ), .A2(\u_ascii_h/_07_ ), .A3(\u_ascii_h/_00_ ), .ZN(\u_ascii_h/_25_ ) );
NAND2_X1 \u_ascii_h/_66_ ( .A1(\u_ascii_h/_13_ ), .A2(\u_ascii_h/_10_ ), .ZN(\u_ascii_h/_26_ ) );
NAND4_X1 \u_ascii_h/_67_ ( .A1(\u_ascii_h/_24_ ), .A2(\u_ascii_h/_04_ ), .A3(\u_ascii_h/_25_ ), .A4(\u_ascii_h/_26_ ), .ZN(\u_ascii_h/_37_ ) );
NAND3_X1 \u_ascii_h/_68_ ( .A1(\u_ascii_h/_10_ ), .A2(\u_ascii_h/_01_ ), .A3(\u_ascii_h/_12_ ), .ZN(\u_ascii_h/_27_ ) );
AOI22_X1 \u_ascii_h/_69_ ( .A1(\u_ascii_h/_08_ ), .A2(\u_ascii_h/_05_ ), .B1(\u_ascii_h/_18_ ), .B2(\u_ascii_h/_21_ ), .ZN(\u_ascii_h/_28_ ) );
NAND4_X1 \u_ascii_h/_70_ ( .A1(\u_ascii_h/_16_ ), .A2(\u_ascii_h/_19_ ), .A3(\u_ascii_h/_27_ ), .A4(\u_ascii_h/_28_ ), .ZN(\u_ascii_h/_38_ ) );
OAI21_X1 \u_ascii_h/_71_ ( .A(\u_ascii_h/_21_ ), .B1(\u_ascii_h/_01_ ), .B2(\u_ascii_h/_12_ ), .ZN(\u_ascii_h/_29_ ) );
NAND3_X1 \u_ascii_h/_72_ ( .A1(\u_ascii_h/_14_ ), .A2(\u_ascii_h/_01_ ), .A3(\u_ascii_h/_12_ ), .ZN(\u_ascii_h/_30_ ) );
NAND3_X1 \u_ascii_h/_73_ ( .A1(\u_ascii_h/_29_ ), .A2(\u_ascii_h/_30_ ), .A3(\u_ascii_h/_04_ ), .ZN(\u_ascii_h/_39_ ) );
AND2_X1 \u_ascii_h/_74_ ( .A1(\u_ascii_h/_12_ ), .A2(\u_ascii_h/_01_ ), .ZN(\u_ascii_h/_31_ ) );
OAI21_X1 \u_ascii_h/_75_ ( .A(\u_ascii_h/_08_ ), .B1(\u_ascii_h/_31_ ), .B2(\u_ascii_h/_13_ ), .ZN(\u_ascii_h/_32_ ) );
NAND2_X1 \u_ascii_h/_76_ ( .A1(\u_ascii_h/_10_ ), .A2(\u_ascii_h/_18_ ), .ZN(\u_ascii_h/_33_ ) );
NAND4_X1 \u_ascii_h/_77_ ( .A1(\u_ascii_h/_32_ ), .A2(\u_ascii_h/_04_ ), .A3(\u_ascii_h/_29_ ), .A4(\u_ascii_h/_33_ ), .ZN(\u_ascii_h/_40_ ) );
AOI22_X1 \u_ascii_h/_78_ ( .A1(\u_ascii_h/_14_ ), .A2(\u_ascii_h/_13_ ), .B1(\u_ascii_h/_08_ ), .B2(\u_ascii_h/_05_ ), .ZN(\u_ascii_h/_34_ ) );
NAND4_X1 \u_ascii_h/_79_ ( .A1(\u_ascii_h/_34_ ), .A2(\u_ascii_h/_04_ ), .A3(\u_ascii_h/_22_ ), .A4(\u_ascii_h/_33_ ), .ZN(\u_ascii_h/_41_ ) );
LOGIC1_X1 \u_ascii_h/_80_ ( .Z(\u_ascii_h/_42_ ) );
BUF_X1 \u_ascii_h/_81_ ( .A(\u_ascii_h/_42_ ), .Z(\ascii_seg [8] ) );
BUF_X1 \u_ascii_h/_82_ ( .A(\ascii_code [7] ), .Z(\u_ascii_h/_03_ ) );
BUF_X1 \u_ascii_h/_83_ ( .A(\ascii_code [6] ), .Z(\u_ascii_h/_02_ ) );
BUF_X1 \u_ascii_h/_84_ ( .A(\ascii_code [5] ), .Z(\u_ascii_h/_01_ ) );
BUF_X1 \u_ascii_h/_85_ ( .A(\ascii_code [4] ), .Z(\u_ascii_h/_00_ ) );
BUF_X1 \u_ascii_h/_86_ ( .A(display_en ), .Z(\u_ascii_h/_04_ ) );
BUF_X1 \u_ascii_h/_87_ ( .A(\u_ascii_h/_35_ ), .Z(\ascii_seg [9] ) );
BUF_X1 \u_ascii_h/_88_ ( .A(\u_ascii_h/_36_ ), .Z(\ascii_seg [10] ) );
BUF_X1 \u_ascii_h/_89_ ( .A(\u_ascii_h/_37_ ), .Z(\ascii_seg [11] ) );
BUF_X1 \u_ascii_h/_90_ ( .A(\u_ascii_h/_38_ ), .Z(\ascii_seg [12] ) );
BUF_X1 \u_ascii_h/_91_ ( .A(\u_ascii_h/_39_ ), .Z(\ascii_seg [13] ) );
BUF_X1 \u_ascii_h/_92_ ( .A(\u_ascii_h/_40_ ), .Z(\ascii_seg [14] ) );
BUF_X1 \u_ascii_h/_93_ ( .A(\u_ascii_h/_41_ ), .Z(\ascii_seg [15] ) );
NOR2_X4 \u_ascii_l/_43_ ( .A1(\u_ascii_l/_01_ ), .A2(\u_ascii_l/_00_ ), .ZN(\u_ascii_l/_05_ ) );
INV_X2 \u_ascii_l/_44_ ( .A(\u_ascii_l/_05_ ), .ZN(\u_ascii_l/_06_ ) );
INV_X4 \u_ascii_l/_45_ ( .A(\u_ascii_l/_02_ ), .ZN(\u_ascii_l/_07_ ) );
NOR2_X2 \u_ascii_l/_46_ ( .A1(\u_ascii_l/_07_ ), .A2(\u_ascii_l/_03_ ), .ZN(\u_ascii_l/_08_ ) );
INV_X16 \u_ascii_l/_47_ ( .A(\u_ascii_l/_03_ ), .ZN(\u_ascii_l/_09_ ) );
NOR2_X2 \u_ascii_l/_48_ ( .A1(\u_ascii_l/_09_ ), .A2(\u_ascii_l/_02_ ), .ZN(\u_ascii_l/_10_ ) );
OR3_X4 \u_ascii_l/_49_ ( .A1(\u_ascii_l/_06_ ), .A2(\u_ascii_l/_08_ ), .A3(\u_ascii_l/_10_ ), .ZN(\u_ascii_l/_11_ ) );
INV_X32 \u_ascii_l/_50_ ( .A(\u_ascii_l/_00_ ), .ZN(\u_ascii_l/_12_ ) );
NOR2_X2 \u_ascii_l/_51_ ( .A1(\u_ascii_l/_12_ ), .A2(\u_ascii_l/_01_ ), .ZN(\u_ascii_l/_13_ ) );
NOR2_X4 \u_ascii_l/_52_ ( .A1(\u_ascii_l/_03_ ), .A2(\u_ascii_l/_02_ ), .ZN(\u_ascii_l/_14_ ) );
AND2_X1 \u_ascii_l/_53_ ( .A1(\u_ascii_l/_13_ ), .A2(\u_ascii_l/_14_ ), .ZN(\u_ascii_l/_15_ ) );
INV_X1 \u_ascii_l/_54_ ( .A(\u_ascii_l/_15_ ), .ZN(\u_ascii_l/_16_ ) );
INV_X1 \u_ascii_l/_55_ ( .A(\u_ascii_l/_04_ ), .ZN(\u_ascii_l/_17_ ) );
AND2_X4 \u_ascii_l/_56_ ( .A1(\u_ascii_l/_01_ ), .A2(\u_ascii_l/_00_ ), .ZN(\u_ascii_l/_18_ ) );
AOI21_X1 \u_ascii_l/_57_ ( .A(\u_ascii_l/_17_ ), .B1(\u_ascii_l/_08_ ), .B2(\u_ascii_l/_18_ ), .ZN(\u_ascii_l/_19_ ) );
NAND3_X1 \u_ascii_l/_58_ ( .A1(\u_ascii_l/_11_ ), .A2(\u_ascii_l/_16_ ), .A3(\u_ascii_l/_19_ ), .ZN(\u_ascii_l/_35_ ) );
NAND2_X1 \u_ascii_l/_59_ ( .A1(\u_ascii_l/_06_ ), .A2(\u_ascii_l/_14_ ), .ZN(\u_ascii_l/_20_ ) );
AND2_X2 \u_ascii_l/_60_ ( .A1(\u_ascii_l/_03_ ), .A2(\u_ascii_l/_02_ ), .ZN(\u_ascii_l/_21_ ) );
NAND2_X1 \u_ascii_l/_61_ ( .A1(\u_ascii_l/_13_ ), .A2(\u_ascii_l/_21_ ), .ZN(\u_ascii_l/_22_ ) );
NAND3_X1 \u_ascii_l/_62_ ( .A1(\u_ascii_l/_19_ ), .A2(\u_ascii_l/_20_ ), .A3(\u_ascii_l/_22_ ), .ZN(\u_ascii_l/_36_ ) );
NOR3_X1 \u_ascii_l/_63_ ( .A1(\u_ascii_l/_07_ ), .A2(\u_ascii_l/_03_ ), .A3(\u_ascii_l/_01_ ), .ZN(\u_ascii_l/_23_ ) );
AOI21_X1 \u_ascii_l/_64_ ( .A(\u_ascii_l/_23_ ), .B1(\u_ascii_l/_08_ ), .B2(\u_ascii_l/_18_ ), .ZN(\u_ascii_l/_24_ ) );
NAND3_X1 \u_ascii_l/_65_ ( .A1(\u_ascii_l/_09_ ), .A2(\u_ascii_l/_07_ ), .A3(\u_ascii_l/_00_ ), .ZN(\u_ascii_l/_25_ ) );
NAND2_X1 \u_ascii_l/_66_ ( .A1(\u_ascii_l/_13_ ), .A2(\u_ascii_l/_10_ ), .ZN(\u_ascii_l/_26_ ) );
NAND4_X1 \u_ascii_l/_67_ ( .A1(\u_ascii_l/_24_ ), .A2(\u_ascii_l/_04_ ), .A3(\u_ascii_l/_25_ ), .A4(\u_ascii_l/_26_ ), .ZN(\u_ascii_l/_37_ ) );
NAND3_X1 \u_ascii_l/_68_ ( .A1(\u_ascii_l/_10_ ), .A2(\u_ascii_l/_01_ ), .A3(\u_ascii_l/_12_ ), .ZN(\u_ascii_l/_27_ ) );
AOI22_X1 \u_ascii_l/_69_ ( .A1(\u_ascii_l/_08_ ), .A2(\u_ascii_l/_05_ ), .B1(\u_ascii_l/_18_ ), .B2(\u_ascii_l/_21_ ), .ZN(\u_ascii_l/_28_ ) );
NAND4_X1 \u_ascii_l/_70_ ( .A1(\u_ascii_l/_16_ ), .A2(\u_ascii_l/_19_ ), .A3(\u_ascii_l/_27_ ), .A4(\u_ascii_l/_28_ ), .ZN(\u_ascii_l/_38_ ) );
OAI21_X1 \u_ascii_l/_71_ ( .A(\u_ascii_l/_21_ ), .B1(\u_ascii_l/_01_ ), .B2(\u_ascii_l/_12_ ), .ZN(\u_ascii_l/_29_ ) );
NAND3_X1 \u_ascii_l/_72_ ( .A1(\u_ascii_l/_14_ ), .A2(\u_ascii_l/_01_ ), .A3(\u_ascii_l/_12_ ), .ZN(\u_ascii_l/_30_ ) );
NAND3_X1 \u_ascii_l/_73_ ( .A1(\u_ascii_l/_29_ ), .A2(\u_ascii_l/_30_ ), .A3(\u_ascii_l/_04_ ), .ZN(\u_ascii_l/_39_ ) );
AND2_X1 \u_ascii_l/_74_ ( .A1(\u_ascii_l/_12_ ), .A2(\u_ascii_l/_01_ ), .ZN(\u_ascii_l/_31_ ) );
OAI21_X1 \u_ascii_l/_75_ ( .A(\u_ascii_l/_08_ ), .B1(\u_ascii_l/_31_ ), .B2(\u_ascii_l/_13_ ), .ZN(\u_ascii_l/_32_ ) );
NAND2_X1 \u_ascii_l/_76_ ( .A1(\u_ascii_l/_10_ ), .A2(\u_ascii_l/_18_ ), .ZN(\u_ascii_l/_33_ ) );
NAND4_X1 \u_ascii_l/_77_ ( .A1(\u_ascii_l/_32_ ), .A2(\u_ascii_l/_04_ ), .A3(\u_ascii_l/_29_ ), .A4(\u_ascii_l/_33_ ), .ZN(\u_ascii_l/_40_ ) );
AOI22_X1 \u_ascii_l/_78_ ( .A1(\u_ascii_l/_14_ ), .A2(\u_ascii_l/_13_ ), .B1(\u_ascii_l/_08_ ), .B2(\u_ascii_l/_05_ ), .ZN(\u_ascii_l/_34_ ) );
NAND4_X1 \u_ascii_l/_79_ ( .A1(\u_ascii_l/_34_ ), .A2(\u_ascii_l/_04_ ), .A3(\u_ascii_l/_22_ ), .A4(\u_ascii_l/_33_ ), .ZN(\u_ascii_l/_41_ ) );
LOGIC1_X1 \u_ascii_l/_80_ ( .Z(\u_ascii_l/_42_ ) );
BUF_X1 \u_ascii_l/_81_ ( .A(\u_ascii_l/_42_ ), .Z(\ascii_seg [0] ) );
BUF_X1 \u_ascii_l/_82_ ( .A(\ascii_code [3] ), .Z(\u_ascii_l/_03_ ) );
BUF_X1 \u_ascii_l/_83_ ( .A(\ascii_code [2] ), .Z(\u_ascii_l/_02_ ) );
BUF_X1 \u_ascii_l/_84_ ( .A(\ascii_code [1] ), .Z(\u_ascii_l/_01_ ) );
BUF_X1 \u_ascii_l/_85_ ( .A(\ascii_code [0] ), .Z(\u_ascii_l/_00_ ) );
BUF_X1 \u_ascii_l/_86_ ( .A(display_en ), .Z(\u_ascii_l/_04_ ) );
BUF_X1 \u_ascii_l/_87_ ( .A(\u_ascii_l/_35_ ), .Z(\ascii_seg [1] ) );
BUF_X1 \u_ascii_l/_88_ ( .A(\u_ascii_l/_36_ ), .Z(\ascii_seg [2] ) );
BUF_X1 \u_ascii_l/_89_ ( .A(\u_ascii_l/_37_ ), .Z(\ascii_seg [3] ) );
BUF_X1 \u_ascii_l/_90_ ( .A(\u_ascii_l/_38_ ), .Z(\ascii_seg [4] ) );
BUF_X1 \u_ascii_l/_91_ ( .A(\u_ascii_l/_39_ ), .Z(\ascii_seg [5] ) );
BUF_X1 \u_ascii_l/_92_ ( .A(\u_ascii_l/_40_ ), .Z(\ascii_seg [6] ) );
BUF_X1 \u_ascii_l/_93_ ( .A(\u_ascii_l/_41_ ), .Z(\ascii_seg [7] ) );
NOR2_X4 \u_count_h/_43_ ( .A1(\u_count_h/_01_ ), .A2(\u_count_h/_00_ ), .ZN(\u_count_h/_05_ ) );
INV_X2 \u_count_h/_44_ ( .A(\u_count_h/_05_ ), .ZN(\u_count_h/_06_ ) );
INV_X4 \u_count_h/_45_ ( .A(\u_count_h/_02_ ), .ZN(\u_count_h/_07_ ) );
NOR2_X2 \u_count_h/_46_ ( .A1(\u_count_h/_07_ ), .A2(\u_count_h/_03_ ), .ZN(\u_count_h/_08_ ) );
INV_X16 \u_count_h/_47_ ( .A(\u_count_h/_03_ ), .ZN(\u_count_h/_09_ ) );
NOR2_X2 \u_count_h/_48_ ( .A1(\u_count_h/_09_ ), .A2(\u_count_h/_02_ ), .ZN(\u_count_h/_10_ ) );
OR3_X4 \u_count_h/_49_ ( .A1(\u_count_h/_06_ ), .A2(\u_count_h/_08_ ), .A3(\u_count_h/_10_ ), .ZN(\u_count_h/_11_ ) );
INV_X32 \u_count_h/_50_ ( .A(\u_count_h/_00_ ), .ZN(\u_count_h/_12_ ) );
NOR2_X2 \u_count_h/_51_ ( .A1(\u_count_h/_12_ ), .A2(\u_count_h/_01_ ), .ZN(\u_count_h/_13_ ) );
NOR2_X4 \u_count_h/_52_ ( .A1(\u_count_h/_03_ ), .A2(\u_count_h/_02_ ), .ZN(\u_count_h/_14_ ) );
AND2_X1 \u_count_h/_53_ ( .A1(\u_count_h/_13_ ), .A2(\u_count_h/_14_ ), .ZN(\u_count_h/_15_ ) );
INV_X1 \u_count_h/_54_ ( .A(\u_count_h/_15_ ), .ZN(\u_count_h/_16_ ) );
INV_X1 \u_count_h/_55_ ( .A(\u_count_h/_04_ ), .ZN(\u_count_h/_17_ ) );
AND2_X4 \u_count_h/_56_ ( .A1(\u_count_h/_01_ ), .A2(\u_count_h/_00_ ), .ZN(\u_count_h/_18_ ) );
AOI21_X1 \u_count_h/_57_ ( .A(\u_count_h/_17_ ), .B1(\u_count_h/_08_ ), .B2(\u_count_h/_18_ ), .ZN(\u_count_h/_19_ ) );
NAND3_X1 \u_count_h/_58_ ( .A1(\u_count_h/_11_ ), .A2(\u_count_h/_16_ ), .A3(\u_count_h/_19_ ), .ZN(\u_count_h/_35_ ) );
NAND2_X1 \u_count_h/_59_ ( .A1(\u_count_h/_06_ ), .A2(\u_count_h/_14_ ), .ZN(\u_count_h/_20_ ) );
AND2_X2 \u_count_h/_60_ ( .A1(\u_count_h/_03_ ), .A2(\u_count_h/_02_ ), .ZN(\u_count_h/_21_ ) );
NAND2_X1 \u_count_h/_61_ ( .A1(\u_count_h/_13_ ), .A2(\u_count_h/_21_ ), .ZN(\u_count_h/_22_ ) );
NAND3_X1 \u_count_h/_62_ ( .A1(\u_count_h/_19_ ), .A2(\u_count_h/_20_ ), .A3(\u_count_h/_22_ ), .ZN(\u_count_h/_36_ ) );
NOR3_X1 \u_count_h/_63_ ( .A1(\u_count_h/_07_ ), .A2(\u_count_h/_03_ ), .A3(\u_count_h/_01_ ), .ZN(\u_count_h/_23_ ) );
AOI21_X1 \u_count_h/_64_ ( .A(\u_count_h/_23_ ), .B1(\u_count_h/_08_ ), .B2(\u_count_h/_18_ ), .ZN(\u_count_h/_24_ ) );
NAND3_X1 \u_count_h/_65_ ( .A1(\u_count_h/_09_ ), .A2(\u_count_h/_07_ ), .A3(\u_count_h/_00_ ), .ZN(\u_count_h/_25_ ) );
NAND2_X1 \u_count_h/_66_ ( .A1(\u_count_h/_13_ ), .A2(\u_count_h/_10_ ), .ZN(\u_count_h/_26_ ) );
NAND4_X1 \u_count_h/_67_ ( .A1(\u_count_h/_24_ ), .A2(\u_count_h/_04_ ), .A3(\u_count_h/_25_ ), .A4(\u_count_h/_26_ ), .ZN(\u_count_h/_37_ ) );
NAND3_X1 \u_count_h/_68_ ( .A1(\u_count_h/_10_ ), .A2(\u_count_h/_01_ ), .A3(\u_count_h/_12_ ), .ZN(\u_count_h/_27_ ) );
AOI22_X1 \u_count_h/_69_ ( .A1(\u_count_h/_08_ ), .A2(\u_count_h/_05_ ), .B1(\u_count_h/_18_ ), .B2(\u_count_h/_21_ ), .ZN(\u_count_h/_28_ ) );
NAND4_X1 \u_count_h/_70_ ( .A1(\u_count_h/_16_ ), .A2(\u_count_h/_19_ ), .A3(\u_count_h/_27_ ), .A4(\u_count_h/_28_ ), .ZN(\u_count_h/_38_ ) );
OAI21_X1 \u_count_h/_71_ ( .A(\u_count_h/_21_ ), .B1(\u_count_h/_01_ ), .B2(\u_count_h/_12_ ), .ZN(\u_count_h/_29_ ) );
NAND3_X1 \u_count_h/_72_ ( .A1(\u_count_h/_14_ ), .A2(\u_count_h/_01_ ), .A3(\u_count_h/_12_ ), .ZN(\u_count_h/_30_ ) );
NAND3_X1 \u_count_h/_73_ ( .A1(\u_count_h/_29_ ), .A2(\u_count_h/_30_ ), .A3(\u_count_h/_04_ ), .ZN(\u_count_h/_39_ ) );
AND2_X1 \u_count_h/_74_ ( .A1(\u_count_h/_12_ ), .A2(\u_count_h/_01_ ), .ZN(\u_count_h/_31_ ) );
OAI21_X1 \u_count_h/_75_ ( .A(\u_count_h/_08_ ), .B1(\u_count_h/_31_ ), .B2(\u_count_h/_13_ ), .ZN(\u_count_h/_32_ ) );
NAND2_X1 \u_count_h/_76_ ( .A1(\u_count_h/_10_ ), .A2(\u_count_h/_18_ ), .ZN(\u_count_h/_33_ ) );
NAND4_X1 \u_count_h/_77_ ( .A1(\u_count_h/_32_ ), .A2(\u_count_h/_04_ ), .A3(\u_count_h/_29_ ), .A4(\u_count_h/_33_ ), .ZN(\u_count_h/_40_ ) );
AOI22_X1 \u_count_h/_78_ ( .A1(\u_count_h/_14_ ), .A2(\u_count_h/_13_ ), .B1(\u_count_h/_08_ ), .B2(\u_count_h/_05_ ), .ZN(\u_count_h/_34_ ) );
NAND4_X1 \u_count_h/_79_ ( .A1(\u_count_h/_34_ ), .A2(\u_count_h/_04_ ), .A3(\u_count_h/_22_ ), .A4(\u_count_h/_33_ ), .ZN(\u_count_h/_41_ ) );
LOGIC1_X1 \u_count_h/_80_ ( .Z(\u_count_h/_42_ ) );
BUF_X1 \u_count_h/_81_ ( .A(\u_count_h/_42_ ), .Z(\count_seg [8] ) );
BUF_X1 \u_count_h/_82_ ( .A(\count [7] ), .Z(\u_count_h/_03_ ) );
BUF_X1 \u_count_h/_83_ ( .A(\count [6] ), .Z(\u_count_h/_02_ ) );
BUF_X1 \u_count_h/_84_ ( .A(\count [5] ), .Z(\u_count_h/_01_ ) );
BUF_X1 \u_count_h/_85_ ( .A(\count [4] ), .Z(\u_count_h/_00_ ) );
BUF_X1 \u_count_h/_86_ ( .A(_141_ ), .Z(\u_count_h/_04_ ) );
BUF_X1 \u_count_h/_87_ ( .A(\u_count_h/_35_ ), .Z(\count_seg [9] ) );
BUF_X1 \u_count_h/_88_ ( .A(\u_count_h/_36_ ), .Z(\count_seg [10] ) );
BUF_X1 \u_count_h/_89_ ( .A(\u_count_h/_37_ ), .Z(\count_seg [11] ) );
BUF_X1 \u_count_h/_90_ ( .A(\u_count_h/_38_ ), .Z(\count_seg [12] ) );
BUF_X1 \u_count_h/_91_ ( .A(\u_count_h/_39_ ), .Z(\count_seg [13] ) );
BUF_X1 \u_count_h/_92_ ( .A(\u_count_h/_40_ ), .Z(\count_seg [14] ) );
BUF_X1 \u_count_h/_93_ ( .A(\u_count_h/_41_ ), .Z(\count_seg [15] ) );
NOR2_X4 \u_count_l/_43_ ( .A1(\u_count_l/_01_ ), .A2(\u_count_l/_00_ ), .ZN(\u_count_l/_05_ ) );
INV_X2 \u_count_l/_44_ ( .A(\u_count_l/_05_ ), .ZN(\u_count_l/_06_ ) );
INV_X4 \u_count_l/_45_ ( .A(\u_count_l/_02_ ), .ZN(\u_count_l/_07_ ) );
NOR2_X2 \u_count_l/_46_ ( .A1(\u_count_l/_07_ ), .A2(\u_count_l/_03_ ), .ZN(\u_count_l/_08_ ) );
INV_X16 \u_count_l/_47_ ( .A(\u_count_l/_03_ ), .ZN(\u_count_l/_09_ ) );
NOR2_X2 \u_count_l/_48_ ( .A1(\u_count_l/_09_ ), .A2(\u_count_l/_02_ ), .ZN(\u_count_l/_10_ ) );
OR3_X4 \u_count_l/_49_ ( .A1(\u_count_l/_06_ ), .A2(\u_count_l/_08_ ), .A3(\u_count_l/_10_ ), .ZN(\u_count_l/_11_ ) );
INV_X32 \u_count_l/_50_ ( .A(\u_count_l/_00_ ), .ZN(\u_count_l/_12_ ) );
NOR2_X2 \u_count_l/_51_ ( .A1(\u_count_l/_12_ ), .A2(\u_count_l/_01_ ), .ZN(\u_count_l/_13_ ) );
NOR2_X4 \u_count_l/_52_ ( .A1(\u_count_l/_03_ ), .A2(\u_count_l/_02_ ), .ZN(\u_count_l/_14_ ) );
AND2_X1 \u_count_l/_53_ ( .A1(\u_count_l/_13_ ), .A2(\u_count_l/_14_ ), .ZN(\u_count_l/_15_ ) );
INV_X1 \u_count_l/_54_ ( .A(\u_count_l/_15_ ), .ZN(\u_count_l/_16_ ) );
INV_X1 \u_count_l/_55_ ( .A(\u_count_l/_04_ ), .ZN(\u_count_l/_17_ ) );
AND2_X4 \u_count_l/_56_ ( .A1(\u_count_l/_01_ ), .A2(\u_count_l/_00_ ), .ZN(\u_count_l/_18_ ) );
AOI21_X1 \u_count_l/_57_ ( .A(\u_count_l/_17_ ), .B1(\u_count_l/_08_ ), .B2(\u_count_l/_18_ ), .ZN(\u_count_l/_19_ ) );
NAND3_X1 \u_count_l/_58_ ( .A1(\u_count_l/_11_ ), .A2(\u_count_l/_16_ ), .A3(\u_count_l/_19_ ), .ZN(\u_count_l/_35_ ) );
NAND2_X1 \u_count_l/_59_ ( .A1(\u_count_l/_06_ ), .A2(\u_count_l/_14_ ), .ZN(\u_count_l/_20_ ) );
AND2_X2 \u_count_l/_60_ ( .A1(\u_count_l/_03_ ), .A2(\u_count_l/_02_ ), .ZN(\u_count_l/_21_ ) );
NAND2_X1 \u_count_l/_61_ ( .A1(\u_count_l/_13_ ), .A2(\u_count_l/_21_ ), .ZN(\u_count_l/_22_ ) );
NAND3_X1 \u_count_l/_62_ ( .A1(\u_count_l/_19_ ), .A2(\u_count_l/_20_ ), .A3(\u_count_l/_22_ ), .ZN(\u_count_l/_36_ ) );
NOR3_X1 \u_count_l/_63_ ( .A1(\u_count_l/_07_ ), .A2(\u_count_l/_03_ ), .A3(\u_count_l/_01_ ), .ZN(\u_count_l/_23_ ) );
AOI21_X1 \u_count_l/_64_ ( .A(\u_count_l/_23_ ), .B1(\u_count_l/_08_ ), .B2(\u_count_l/_18_ ), .ZN(\u_count_l/_24_ ) );
NAND3_X1 \u_count_l/_65_ ( .A1(\u_count_l/_09_ ), .A2(\u_count_l/_07_ ), .A3(\u_count_l/_00_ ), .ZN(\u_count_l/_25_ ) );
NAND2_X1 \u_count_l/_66_ ( .A1(\u_count_l/_13_ ), .A2(\u_count_l/_10_ ), .ZN(\u_count_l/_26_ ) );
NAND4_X1 \u_count_l/_67_ ( .A1(\u_count_l/_24_ ), .A2(\u_count_l/_04_ ), .A3(\u_count_l/_25_ ), .A4(\u_count_l/_26_ ), .ZN(\u_count_l/_37_ ) );
NAND3_X1 \u_count_l/_68_ ( .A1(\u_count_l/_10_ ), .A2(\u_count_l/_01_ ), .A3(\u_count_l/_12_ ), .ZN(\u_count_l/_27_ ) );
AOI22_X1 \u_count_l/_69_ ( .A1(\u_count_l/_08_ ), .A2(\u_count_l/_05_ ), .B1(\u_count_l/_18_ ), .B2(\u_count_l/_21_ ), .ZN(\u_count_l/_28_ ) );
NAND4_X1 \u_count_l/_70_ ( .A1(\u_count_l/_16_ ), .A2(\u_count_l/_19_ ), .A3(\u_count_l/_27_ ), .A4(\u_count_l/_28_ ), .ZN(\u_count_l/_38_ ) );
OAI21_X1 \u_count_l/_71_ ( .A(\u_count_l/_21_ ), .B1(\u_count_l/_01_ ), .B2(\u_count_l/_12_ ), .ZN(\u_count_l/_29_ ) );
NAND3_X1 \u_count_l/_72_ ( .A1(\u_count_l/_14_ ), .A2(\u_count_l/_01_ ), .A3(\u_count_l/_12_ ), .ZN(\u_count_l/_30_ ) );
NAND3_X1 \u_count_l/_73_ ( .A1(\u_count_l/_29_ ), .A2(\u_count_l/_30_ ), .A3(\u_count_l/_04_ ), .ZN(\u_count_l/_39_ ) );
AND2_X1 \u_count_l/_74_ ( .A1(\u_count_l/_12_ ), .A2(\u_count_l/_01_ ), .ZN(\u_count_l/_31_ ) );
OAI21_X1 \u_count_l/_75_ ( .A(\u_count_l/_08_ ), .B1(\u_count_l/_31_ ), .B2(\u_count_l/_13_ ), .ZN(\u_count_l/_32_ ) );
NAND2_X1 \u_count_l/_76_ ( .A1(\u_count_l/_10_ ), .A2(\u_count_l/_18_ ), .ZN(\u_count_l/_33_ ) );
NAND4_X1 \u_count_l/_77_ ( .A1(\u_count_l/_32_ ), .A2(\u_count_l/_04_ ), .A3(\u_count_l/_29_ ), .A4(\u_count_l/_33_ ), .ZN(\u_count_l/_40_ ) );
AOI22_X1 \u_count_l/_78_ ( .A1(\u_count_l/_14_ ), .A2(\u_count_l/_13_ ), .B1(\u_count_l/_08_ ), .B2(\u_count_l/_05_ ), .ZN(\u_count_l/_34_ ) );
NAND4_X1 \u_count_l/_79_ ( .A1(\u_count_l/_34_ ), .A2(\u_count_l/_04_ ), .A3(\u_count_l/_22_ ), .A4(\u_count_l/_33_ ), .ZN(\u_count_l/_41_ ) );
LOGIC1_X1 \u_count_l/_80_ ( .Z(\u_count_l/_42_ ) );
BUF_X1 \u_count_l/_81_ ( .A(\u_count_l/_42_ ), .Z(\count_seg [0] ) );
BUF_X1 \u_count_l/_82_ ( .A(\count [3] ), .Z(\u_count_l/_03_ ) );
BUF_X1 \u_count_l/_83_ ( .A(\count [2] ), .Z(\u_count_l/_02_ ) );
BUF_X1 \u_count_l/_84_ ( .A(\count [1] ), .Z(\u_count_l/_01_ ) );
BUF_X1 \u_count_l/_85_ ( .A(\count [0] ), .Z(\u_count_l/_00_ ) );
BUF_X1 \u_count_l/_86_ ( .A(_141_ ), .Z(\u_count_l/_04_ ) );
BUF_X1 \u_count_l/_87_ ( .A(\u_count_l/_35_ ), .Z(\count_seg [1] ) );
BUF_X1 \u_count_l/_88_ ( .A(\u_count_l/_36_ ), .Z(\count_seg [2] ) );
BUF_X1 \u_count_l/_89_ ( .A(\u_count_l/_37_ ), .Z(\count_seg [3] ) );
BUF_X1 \u_count_l/_90_ ( .A(\u_count_l/_38_ ), .Z(\count_seg [4] ) );
BUF_X1 \u_count_l/_91_ ( .A(\u_count_l/_39_ ), .Z(\count_seg [5] ) );
BUF_X1 \u_count_l/_92_ ( .A(\u_count_l/_40_ ), .Z(\count_seg [6] ) );
BUF_X1 \u_count_l/_93_ ( .A(\u_count_l/_41_ ), .Z(\count_seg [7] ) );
MUX2_X1 \u_ps2_keyboard/_0528_ ( .A(\u_ps2_keyboard/_0222_ ), .B(\u_ps2_keyboard/_0230_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0270_ ) );
MUX2_X1 \u_ps2_keyboard/_0529_ ( .A(\u_ps2_keyboard/_0206_ ), .B(\u_ps2_keyboard/_0214_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0271_ ) );
INV_X2 \u_ps2_keyboard/_0530_ ( .A(\u_ps2_keyboard/_0434_ ), .ZN(\u_ps2_keyboard/_0272_ ) );
MUX2_X1 \u_ps2_keyboard/_0531_ ( .A(\u_ps2_keyboard/_0270_ ), .B(\u_ps2_keyboard/_0271_ ), .S(\u_ps2_keyboard/_0272_ ), .Z(\u_ps2_keyboard/_0273_ ) );
MUX2_X1 \u_ps2_keyboard/_0532_ ( .A(\u_ps2_keyboard/_0238_ ), .B(\u_ps2_keyboard/_0254_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0274_ ) );
MUX2_X1 \u_ps2_keyboard/_0533_ ( .A(\u_ps2_keyboard/_0246_ ), .B(\u_ps2_keyboard/_0262_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0275_ ) );
MUX2_X1 \u_ps2_keyboard/_0534_ ( .A(\u_ps2_keyboard/_0274_ ), .B(\u_ps2_keyboard/_0275_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0276_ ) );
MUX2_X1 \u_ps2_keyboard/_0535_ ( .A(\u_ps2_keyboard/_0273_ ), .B(\u_ps2_keyboard/_0276_ ), .S(\u_ps2_keyboard/_0435_ ), .Z(\u_ps2_keyboard/_0438_ ) );
MUX2_X1 \u_ps2_keyboard/_0536_ ( .A(\u_ps2_keyboard/_0223_ ), .B(\u_ps2_keyboard/_0231_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0277_ ) );
MUX2_X1 \u_ps2_keyboard/_0537_ ( .A(\u_ps2_keyboard/_0207_ ), .B(\u_ps2_keyboard/_0215_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0278_ ) );
MUX2_X1 \u_ps2_keyboard/_0538_ ( .A(\u_ps2_keyboard/_0277_ ), .B(\u_ps2_keyboard/_0278_ ), .S(\u_ps2_keyboard/_0272_ ), .Z(\u_ps2_keyboard/_0279_ ) );
MUX2_X1 \u_ps2_keyboard/_0539_ ( .A(\u_ps2_keyboard/_0239_ ), .B(\u_ps2_keyboard/_0255_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0280_ ) );
MUX2_X1 \u_ps2_keyboard/_0540_ ( .A(\u_ps2_keyboard/_0247_ ), .B(\u_ps2_keyboard/_0263_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0281_ ) );
MUX2_X1 \u_ps2_keyboard/_0541_ ( .A(\u_ps2_keyboard/_0280_ ), .B(\u_ps2_keyboard/_0281_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0282_ ) );
MUX2_X1 \u_ps2_keyboard/_0542_ ( .A(\u_ps2_keyboard/_0279_ ), .B(\u_ps2_keyboard/_0282_ ), .S(\u_ps2_keyboard/_0435_ ), .Z(\u_ps2_keyboard/_0439_ ) );
MUX2_X1 \u_ps2_keyboard/_0543_ ( .A(\u_ps2_keyboard/_0224_ ), .B(\u_ps2_keyboard/_0232_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0283_ ) );
MUX2_X1 \u_ps2_keyboard/_0544_ ( .A(\u_ps2_keyboard/_0208_ ), .B(\u_ps2_keyboard/_0216_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0284_ ) );
MUX2_X1 \u_ps2_keyboard/_0545_ ( .A(\u_ps2_keyboard/_0283_ ), .B(\u_ps2_keyboard/_0284_ ), .S(\u_ps2_keyboard/_0272_ ), .Z(\u_ps2_keyboard/_0285_ ) );
MUX2_X1 \u_ps2_keyboard/_0546_ ( .A(\u_ps2_keyboard/_0240_ ), .B(\u_ps2_keyboard/_0256_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0286_ ) );
MUX2_X1 \u_ps2_keyboard/_0547_ ( .A(\u_ps2_keyboard/_0248_ ), .B(\u_ps2_keyboard/_0264_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0287_ ) );
MUX2_X1 \u_ps2_keyboard/_0548_ ( .A(\u_ps2_keyboard/_0286_ ), .B(\u_ps2_keyboard/_0287_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0288_ ) );
MUX2_X1 \u_ps2_keyboard/_0549_ ( .A(\u_ps2_keyboard/_0285_ ), .B(\u_ps2_keyboard/_0288_ ), .S(\u_ps2_keyboard/_0435_ ), .Z(\u_ps2_keyboard/_0440_ ) );
MUX2_X1 \u_ps2_keyboard/_0550_ ( .A(\u_ps2_keyboard/_0225_ ), .B(\u_ps2_keyboard/_0233_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0289_ ) );
MUX2_X1 \u_ps2_keyboard/_0551_ ( .A(\u_ps2_keyboard/_0209_ ), .B(\u_ps2_keyboard/_0217_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0290_ ) );
MUX2_X1 \u_ps2_keyboard/_0552_ ( .A(\u_ps2_keyboard/_0289_ ), .B(\u_ps2_keyboard/_0290_ ), .S(\u_ps2_keyboard/_0272_ ), .Z(\u_ps2_keyboard/_0291_ ) );
MUX2_X1 \u_ps2_keyboard/_0553_ ( .A(\u_ps2_keyboard/_0241_ ), .B(\u_ps2_keyboard/_0257_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0292_ ) );
MUX2_X1 \u_ps2_keyboard/_0554_ ( .A(\u_ps2_keyboard/_0249_ ), .B(\u_ps2_keyboard/_0265_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0293_ ) );
MUX2_X1 \u_ps2_keyboard/_0555_ ( .A(\u_ps2_keyboard/_0292_ ), .B(\u_ps2_keyboard/_0293_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0294_ ) );
MUX2_X1 \u_ps2_keyboard/_0556_ ( .A(\u_ps2_keyboard/_0291_ ), .B(\u_ps2_keyboard/_0294_ ), .S(\u_ps2_keyboard/_0435_ ), .Z(\u_ps2_keyboard/_0441_ ) );
MUX2_X1 \u_ps2_keyboard/_0557_ ( .A(\u_ps2_keyboard/_0226_ ), .B(\u_ps2_keyboard/_0234_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0295_ ) );
MUX2_X1 \u_ps2_keyboard/_0558_ ( .A(\u_ps2_keyboard/_0210_ ), .B(\u_ps2_keyboard/_0218_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0296_ ) );
MUX2_X1 \u_ps2_keyboard/_0559_ ( .A(\u_ps2_keyboard/_0295_ ), .B(\u_ps2_keyboard/_0296_ ), .S(\u_ps2_keyboard/_0272_ ), .Z(\u_ps2_keyboard/_0297_ ) );
MUX2_X1 \u_ps2_keyboard/_0560_ ( .A(\u_ps2_keyboard/_0242_ ), .B(\u_ps2_keyboard/_0258_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0298_ ) );
MUX2_X1 \u_ps2_keyboard/_0561_ ( .A(\u_ps2_keyboard/_0250_ ), .B(\u_ps2_keyboard/_0266_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0299_ ) );
MUX2_X1 \u_ps2_keyboard/_0562_ ( .A(\u_ps2_keyboard/_0298_ ), .B(\u_ps2_keyboard/_0299_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0300_ ) );
MUX2_X1 \u_ps2_keyboard/_0563_ ( .A(\u_ps2_keyboard/_0297_ ), .B(\u_ps2_keyboard/_0300_ ), .S(\u_ps2_keyboard/_0435_ ), .Z(\u_ps2_keyboard/_0442_ ) );
MUX2_X1 \u_ps2_keyboard/_0564_ ( .A(\u_ps2_keyboard/_0227_ ), .B(\u_ps2_keyboard/_0235_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0301_ ) );
MUX2_X1 \u_ps2_keyboard/_0565_ ( .A(\u_ps2_keyboard/_0211_ ), .B(\u_ps2_keyboard/_0219_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0302_ ) );
MUX2_X1 \u_ps2_keyboard/_0566_ ( .A(\u_ps2_keyboard/_0301_ ), .B(\u_ps2_keyboard/_0302_ ), .S(\u_ps2_keyboard/_0272_ ), .Z(\u_ps2_keyboard/_0303_ ) );
MUX2_X1 \u_ps2_keyboard/_0567_ ( .A(\u_ps2_keyboard/_0243_ ), .B(\u_ps2_keyboard/_0259_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0304_ ) );
MUX2_X1 \u_ps2_keyboard/_0568_ ( .A(\u_ps2_keyboard/_0251_ ), .B(\u_ps2_keyboard/_0267_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0305_ ) );
MUX2_X1 \u_ps2_keyboard/_0569_ ( .A(\u_ps2_keyboard/_0304_ ), .B(\u_ps2_keyboard/_0305_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0306_ ) );
MUX2_X1 \u_ps2_keyboard/_0570_ ( .A(\u_ps2_keyboard/_0303_ ), .B(\u_ps2_keyboard/_0306_ ), .S(\u_ps2_keyboard/_0435_ ), .Z(\u_ps2_keyboard/_0443_ ) );
MUX2_X1 \u_ps2_keyboard/_0571_ ( .A(\u_ps2_keyboard/_0228_ ), .B(\u_ps2_keyboard/_0236_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0307_ ) );
MUX2_X1 \u_ps2_keyboard/_0572_ ( .A(\u_ps2_keyboard/_0212_ ), .B(\u_ps2_keyboard/_0220_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0308_ ) );
MUX2_X1 \u_ps2_keyboard/_0573_ ( .A(\u_ps2_keyboard/_0307_ ), .B(\u_ps2_keyboard/_0308_ ), .S(\u_ps2_keyboard/_0272_ ), .Z(\u_ps2_keyboard/_0309_ ) );
MUX2_X1 \u_ps2_keyboard/_0574_ ( .A(\u_ps2_keyboard/_0244_ ), .B(\u_ps2_keyboard/_0260_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0310_ ) );
MUX2_X1 \u_ps2_keyboard/_0575_ ( .A(\u_ps2_keyboard/_0252_ ), .B(\u_ps2_keyboard/_0268_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0311_ ) );
MUX2_X1 \u_ps2_keyboard/_0576_ ( .A(\u_ps2_keyboard/_0310_ ), .B(\u_ps2_keyboard/_0311_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0312_ ) );
MUX2_X1 \u_ps2_keyboard/_0577_ ( .A(\u_ps2_keyboard/_0309_ ), .B(\u_ps2_keyboard/_0312_ ), .S(\u_ps2_keyboard/_0435_ ), .Z(\u_ps2_keyboard/_0444_ ) );
MUX2_X1 \u_ps2_keyboard/_0578_ ( .A(\u_ps2_keyboard/_0229_ ), .B(\u_ps2_keyboard/_0237_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0313_ ) );
MUX2_X1 \u_ps2_keyboard/_0579_ ( .A(\u_ps2_keyboard/_0213_ ), .B(\u_ps2_keyboard/_0221_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0314_ ) );
MUX2_X1 \u_ps2_keyboard/_0580_ ( .A(\u_ps2_keyboard/_0313_ ), .B(\u_ps2_keyboard/_0314_ ), .S(\u_ps2_keyboard/_0272_ ), .Z(\u_ps2_keyboard/_0315_ ) );
MUX2_X1 \u_ps2_keyboard/_0581_ ( .A(\u_ps2_keyboard/_0245_ ), .B(\u_ps2_keyboard/_0261_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0316_ ) );
MUX2_X1 \u_ps2_keyboard/_0582_ ( .A(\u_ps2_keyboard/_0253_ ), .B(\u_ps2_keyboard/_0269_ ), .S(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0317_ ) );
MUX2_X1 \u_ps2_keyboard/_0583_ ( .A(\u_ps2_keyboard/_0316_ ), .B(\u_ps2_keyboard/_0317_ ), .S(\u_ps2_keyboard/_0433_ ), .Z(\u_ps2_keyboard/_0318_ ) );
MUX2_X1 \u_ps2_keyboard/_0584_ ( .A(\u_ps2_keyboard/_0315_ ), .B(\u_ps2_keyboard/_0318_ ), .S(\u_ps2_keyboard/_0435_ ), .Z(\u_ps2_keyboard/_0445_ ) );
INV_X1 \u_ps2_keyboard/_0585_ ( .A(\u_ps2_keyboard/_0431_ ), .ZN(\u_ps2_keyboard/_0319_ ) );
NOR2_X1 \u_ps2_keyboard/_0586_ ( .A1(\u_ps2_keyboard/_0319_ ), .A2(\u_ps2_keyboard/_0430_ ), .ZN(\u_ps2_keyboard/_0320_ ) );
INV_X1 \u_ps2_keyboard/_0587_ ( .A(\u_ps2_keyboard/_0202_ ), .ZN(\u_ps2_keyboard/_0321_ ) );
NOR2_X1 \u_ps2_keyboard/_0588_ ( .A1(\u_ps2_keyboard/_0321_ ), .A2(\u_ps2_keyboard/_0203_ ), .ZN(\u_ps2_keyboard/_0322_ ) );
AND2_X1 \u_ps2_keyboard/_0589_ ( .A1(\u_ps2_keyboard/_0320_ ), .A2(\u_ps2_keyboard/_0322_ ), .ZN(\u_ps2_keyboard/_0323_ ) );
INV_X1 \u_ps2_keyboard/_0590_ ( .A(\u_ps2_keyboard/_0323_ ), .ZN(\u_ps2_keyboard/_0324_ ) );
INV_X1 \u_ps2_keyboard/_0591_ ( .A(\u_ps2_keyboard/_0204_ ), .ZN(\u_ps2_keyboard/_0325_ ) );
NAND3_X1 \u_ps2_keyboard/_0592_ ( .A1(\u_ps2_keyboard/_0325_ ), .A2(\u_ps2_keyboard/_0437_ ), .A3(\u_ps2_keyboard/_0205_ ), .ZN(\u_ps2_keyboard/_0326_ ) );
NOR2_X1 \u_ps2_keyboard/_0593_ ( .A1(\u_ps2_keyboard/_0324_ ), .A2(\u_ps2_keyboard/_0326_ ), .ZN(\u_ps2_keyboard/_0327_ ) );
MUX2_X1 \u_ps2_keyboard/_0594_ ( .A(\u_ps2_keyboard/_0201_ ), .B(\u_ps2_keyboard/_0432_ ), .S(\u_ps2_keyboard/_0327_ ), .Z(\u_ps2_keyboard/_0105_ ) );
NOR2_X1 \u_ps2_keyboard/_0595_ ( .A1(\u_ps2_keyboard/_0202_ ), .A2(\u_ps2_keyboard/_0203_ ), .ZN(\u_ps2_keyboard/_0328_ ) );
AND2_X1 \u_ps2_keyboard/_0596_ ( .A1(\u_ps2_keyboard/_0320_ ), .A2(\u_ps2_keyboard/_0328_ ), .ZN(\u_ps2_keyboard/_0329_ ) );
INV_X1 \u_ps2_keyboard/_0597_ ( .A(\u_ps2_keyboard/_0329_ ), .ZN(\u_ps2_keyboard/_0330_ ) );
NOR2_X1 \u_ps2_keyboard/_0598_ ( .A1(\u_ps2_keyboard/_0330_ ), .A2(\u_ps2_keyboard/_0326_ ), .ZN(\u_ps2_keyboard/_0331_ ) );
MUX2_X1 \u_ps2_keyboard/_0599_ ( .A(\u_ps2_keyboard/_0200_ ), .B(\u_ps2_keyboard/_0432_ ), .S(\u_ps2_keyboard/_0331_ ), .Z(\u_ps2_keyboard/_0104_ ) );
AND2_X1 \u_ps2_keyboard/_0600_ ( .A1(\u_ps2_keyboard/_0202_ ), .A2(\u_ps2_keyboard/_0203_ ), .ZN(\u_ps2_keyboard/_0332_ ) );
NAND3_X1 \u_ps2_keyboard/_0601_ ( .A1(\u_ps2_keyboard/_0320_ ), .A2(\u_ps2_keyboard/_0204_ ), .A3(\u_ps2_keyboard/_0332_ ), .ZN(\u_ps2_keyboard/_0333_ ) );
INV_X1 \u_ps2_keyboard/_0602_ ( .A(\u_ps2_keyboard/_0205_ ), .ZN(\u_ps2_keyboard/_0334_ ) );
NAND2_X1 \u_ps2_keyboard/_0603_ ( .A1(\u_ps2_keyboard/_0334_ ), .A2(\u_ps2_keyboard/_0437_ ), .ZN(\u_ps2_keyboard/_0335_ ) );
NOR2_X1 \u_ps2_keyboard/_0604_ ( .A1(\u_ps2_keyboard/_0333_ ), .A2(\u_ps2_keyboard/_0335_ ), .ZN(\u_ps2_keyboard/_0336_ ) );
MUX2_X1 \u_ps2_keyboard/_0605_ ( .A(\u_ps2_keyboard/_0199_ ), .B(\u_ps2_keyboard/_0432_ ), .S(\u_ps2_keyboard/_0336_ ), .Z(\u_ps2_keyboard/_0103_ ) );
AND3_X1 \u_ps2_keyboard/_0606_ ( .A1(\u_ps2_keyboard/_0320_ ), .A2(\u_ps2_keyboard/_0321_ ), .A3(\u_ps2_keyboard/_0203_ ), .ZN(\u_ps2_keyboard/_0337_ ) );
NOR2_X1 \u_ps2_keyboard/_0607_ ( .A1(\u_ps2_keyboard/_0335_ ), .A2(\u_ps2_keyboard/_0325_ ), .ZN(\u_ps2_keyboard/_0338_ ) );
NAND2_X1 \u_ps2_keyboard/_0608_ ( .A1(\u_ps2_keyboard/_0337_ ), .A2(\u_ps2_keyboard/_0338_ ), .ZN(\u_ps2_keyboard/_0339_ ) );
MUX2_X1 \u_ps2_keyboard/_0609_ ( .A(\u_ps2_keyboard/_0432_ ), .B(\u_ps2_keyboard/_0198_ ), .S(\u_ps2_keyboard/_0339_ ), .Z(\u_ps2_keyboard/_0102_ ) );
NAND2_X1 \u_ps2_keyboard/_0610_ ( .A1(\u_ps2_keyboard/_0323_ ), .A2(\u_ps2_keyboard/_0338_ ), .ZN(\u_ps2_keyboard/_0340_ ) );
MUX2_X1 \u_ps2_keyboard/_0611_ ( .A(\u_ps2_keyboard/_0432_ ), .B(\u_ps2_keyboard/_0197_ ), .S(\u_ps2_keyboard/_0340_ ), .Z(\u_ps2_keyboard/_0101_ ) );
NAND2_X1 \u_ps2_keyboard/_0612_ ( .A1(\u_ps2_keyboard/_0329_ ), .A2(\u_ps2_keyboard/_0338_ ), .ZN(\u_ps2_keyboard/_0341_ ) );
MUX2_X1 \u_ps2_keyboard/_0613_ ( .A(\u_ps2_keyboard/_0432_ ), .B(\u_ps2_keyboard/_0196_ ), .S(\u_ps2_keyboard/_0341_ ), .Z(\u_ps2_keyboard/_0100_ ) );
INV_X1 \u_ps2_keyboard/_0614_ ( .A(\u_ps2_keyboard/_0432_ ), .ZN(\u_ps2_keyboard/_0342_ ) );
XOR2_X2 \u_ps2_keyboard/_0615_ ( .A(\u_ps2_keyboard/_0193_ ), .B(\u_ps2_keyboard/_0195_ ), .Z(\u_ps2_keyboard/_0343_ ) );
XNOR2_X2 \u_ps2_keyboard/_0616_ ( .A(\u_ps2_keyboard/_0196_ ), .B(\u_ps2_keyboard/_0194_ ), .ZN(\u_ps2_keyboard/_0344_ ) );
XNOR2_X2 \u_ps2_keyboard/_0617_ ( .A(\u_ps2_keyboard/_0343_ ), .B(\u_ps2_keyboard/_0344_ ), .ZN(\u_ps2_keyboard/_0345_ ) );
XNOR2_X1 \u_ps2_keyboard/_0618_ ( .A(\u_ps2_keyboard/_0200_ ), .B(\u_ps2_keyboard/_0199_ ), .ZN(\u_ps2_keyboard/_0346_ ) );
XNOR2_X2 \u_ps2_keyboard/_0619_ ( .A(\u_ps2_keyboard/_0198_ ), .B(\u_ps2_keyboard/_0197_ ), .ZN(\u_ps2_keyboard/_0347_ ) );
XNOR2_X1 \u_ps2_keyboard/_0620_ ( .A(\u_ps2_keyboard/_0346_ ), .B(\u_ps2_keyboard/_0347_ ), .ZN(\u_ps2_keyboard/_0348_ ) );
XNOR2_X2 \u_ps2_keyboard/_0621_ ( .A(\u_ps2_keyboard/_0345_ ), .B(\u_ps2_keyboard/_0348_ ), .ZN(\u_ps2_keyboard/_0349_ ) );
AOI211_X2 \u_ps2_keyboard/_0622_ ( .A(\u_ps2_keyboard/_0342_ ), .B(\u_ps2_keyboard/_0192_ ), .C1(\u_ps2_keyboard/_0349_ ), .C2(\u_ps2_keyboard/_0201_ ), .ZN(\u_ps2_keyboard/_0350_ ) );
OR2_X1 \u_ps2_keyboard/_0623_ ( .A1(\u_ps2_keyboard/_0349_ ), .A2(\u_ps2_keyboard/_0201_ ), .ZN(\u_ps2_keyboard/_0351_ ) );
AND2_X2 \u_ps2_keyboard/_0624_ ( .A1(\u_ps2_keyboard/_0350_ ), .A2(\u_ps2_keyboard/_0351_ ), .ZN(\u_ps2_keyboard/_0352_ ) );
AND2_X1 \u_ps2_keyboard/_0625_ ( .A1(\u_ps2_keyboard/_0321_ ), .A2(\u_ps2_keyboard/_0203_ ), .ZN(\u_ps2_keyboard/_0353_ ) );
NOR2_X1 \u_ps2_keyboard/_0626_ ( .A1(\u_ps2_keyboard/_0334_ ), .A2(\u_ps2_keyboard/_0204_ ), .ZN(\u_ps2_keyboard/_0354_ ) );
AND2_X1 \u_ps2_keyboard/_0627_ ( .A1(\u_ps2_keyboard/_0353_ ), .A2(\u_ps2_keyboard/_0354_ ), .ZN(\u_ps2_keyboard/_0355_ ) );
AND2_X4 \u_ps2_keyboard/_0628_ ( .A1(\u_ps2_keyboard/_0352_ ), .A2(\u_ps2_keyboard/_0355_ ), .ZN(\u_ps2_keyboard/_0356_ ) );
AND2_X4 \u_ps2_keyboard/_0629_ ( .A1(\u_ps2_keyboard/_0356_ ), .A2(\u_ps2_keyboard/_0320_ ), .ZN(\u_ps2_keyboard/_0357_ ) );
NAND2_X4 \u_ps2_keyboard/_0630_ ( .A1(\u_ps2_keyboard/_0357_ ), .A2(\u_ps2_keyboard/_0437_ ), .ZN(\u_ps2_keyboard/_0358_ ) );
NAND3_X1 \u_ps2_keyboard/_0631_ ( .A1(\u_ps2_keyboard/_0448_ ), .A2(\u_ps2_keyboard/_0447_ ), .A3(\u_ps2_keyboard/_0446_ ), .ZN(\u_ps2_keyboard/_0359_ ) );
NOR2_X4 \u_ps2_keyboard/_0632_ ( .A1(\u_ps2_keyboard/_0358_ ), .A2(\u_ps2_keyboard/_0359_ ), .ZN(\u_ps2_keyboard/_0360_ ) );
MUX2_X1 \u_ps2_keyboard/_0633_ ( .A(\u_ps2_keyboard/_0262_ ), .B(\u_ps2_keyboard/_0193_ ), .S(\u_ps2_keyboard/_0360_ ), .Z(\u_ps2_keyboard/_0174_ ) );
MUX2_X1 \u_ps2_keyboard/_0634_ ( .A(\u_ps2_keyboard/_0263_ ), .B(\u_ps2_keyboard/_0194_ ), .S(\u_ps2_keyboard/_0360_ ), .Z(\u_ps2_keyboard/_0175_ ) );
MUX2_X1 \u_ps2_keyboard/_0635_ ( .A(\u_ps2_keyboard/_0264_ ), .B(\u_ps2_keyboard/_0195_ ), .S(\u_ps2_keyboard/_0360_ ), .Z(\u_ps2_keyboard/_0176_ ) );
MUX2_X1 \u_ps2_keyboard/_0636_ ( .A(\u_ps2_keyboard/_0265_ ), .B(\u_ps2_keyboard/_0196_ ), .S(\u_ps2_keyboard/_0360_ ), .Z(\u_ps2_keyboard/_0177_ ) );
MUX2_X1 \u_ps2_keyboard/_0637_ ( .A(\u_ps2_keyboard/_0266_ ), .B(\u_ps2_keyboard/_0197_ ), .S(\u_ps2_keyboard/_0360_ ), .Z(\u_ps2_keyboard/_0178_ ) );
MUX2_X1 \u_ps2_keyboard/_0638_ ( .A(\u_ps2_keyboard/_0267_ ), .B(\u_ps2_keyboard/_0198_ ), .S(\u_ps2_keyboard/_0360_ ), .Z(\u_ps2_keyboard/_0179_ ) );
MUX2_X1 \u_ps2_keyboard/_0639_ ( .A(\u_ps2_keyboard/_0268_ ), .B(\u_ps2_keyboard/_0199_ ), .S(\u_ps2_keyboard/_0360_ ), .Z(\u_ps2_keyboard/_0180_ ) );
MUX2_X1 \u_ps2_keyboard/_0640_ ( .A(\u_ps2_keyboard/_0269_ ), .B(\u_ps2_keyboard/_0200_ ), .S(\u_ps2_keyboard/_0360_ ), .Z(\u_ps2_keyboard/_0181_ ) );
NOR2_X1 \u_ps2_keyboard/_0641_ ( .A1(\u_ps2_keyboard/_0335_ ), .A2(\u_ps2_keyboard/_0204_ ), .ZN(\u_ps2_keyboard/_0361_ ) );
NAND3_X1 \u_ps2_keyboard/_0642_ ( .A1(\u_ps2_keyboard/_0361_ ), .A2(\u_ps2_keyboard/_0320_ ), .A3(\u_ps2_keyboard/_0332_ ), .ZN(\u_ps2_keyboard/_0362_ ) );
MUX2_X1 \u_ps2_keyboard/_0643_ ( .A(\u_ps2_keyboard/_0432_ ), .B(\u_ps2_keyboard/_0195_ ), .S(\u_ps2_keyboard/_0362_ ), .Z(\u_ps2_keyboard/_0099_ ) );
INV_X1 \u_ps2_keyboard/_0644_ ( .A(\u_ps2_keyboard/_0446_ ), .ZN(\u_ps2_keyboard/_0363_ ) );
NAND3_X1 \u_ps2_keyboard/_0645_ ( .A1(\u_ps2_keyboard/_0363_ ), .A2(\u_ps2_keyboard/_0448_ ), .A3(\u_ps2_keyboard/_0447_ ), .ZN(\u_ps2_keyboard/_0364_ ) );
NOR2_X4 \u_ps2_keyboard/_0646_ ( .A1(\u_ps2_keyboard/_0358_ ), .A2(\u_ps2_keyboard/_0364_ ), .ZN(\u_ps2_keyboard/_0365_ ) );
MUX2_X1 \u_ps2_keyboard/_0647_ ( .A(\u_ps2_keyboard/_0254_ ), .B(\u_ps2_keyboard/_0193_ ), .S(\u_ps2_keyboard/_0365_ ), .Z(\u_ps2_keyboard/_0166_ ) );
MUX2_X1 \u_ps2_keyboard/_0648_ ( .A(\u_ps2_keyboard/_0255_ ), .B(\u_ps2_keyboard/_0194_ ), .S(\u_ps2_keyboard/_0365_ ), .Z(\u_ps2_keyboard/_0167_ ) );
MUX2_X1 \u_ps2_keyboard/_0649_ ( .A(\u_ps2_keyboard/_0256_ ), .B(\u_ps2_keyboard/_0195_ ), .S(\u_ps2_keyboard/_0365_ ), .Z(\u_ps2_keyboard/_0168_ ) );
MUX2_X1 \u_ps2_keyboard/_0650_ ( .A(\u_ps2_keyboard/_0257_ ), .B(\u_ps2_keyboard/_0196_ ), .S(\u_ps2_keyboard/_0365_ ), .Z(\u_ps2_keyboard/_0169_ ) );
MUX2_X1 \u_ps2_keyboard/_0651_ ( .A(\u_ps2_keyboard/_0258_ ), .B(\u_ps2_keyboard/_0197_ ), .S(\u_ps2_keyboard/_0365_ ), .Z(\u_ps2_keyboard/_0170_ ) );
MUX2_X1 \u_ps2_keyboard/_0652_ ( .A(\u_ps2_keyboard/_0259_ ), .B(\u_ps2_keyboard/_0198_ ), .S(\u_ps2_keyboard/_0365_ ), .Z(\u_ps2_keyboard/_0171_ ) );
MUX2_X1 \u_ps2_keyboard/_0653_ ( .A(\u_ps2_keyboard/_0260_ ), .B(\u_ps2_keyboard/_0199_ ), .S(\u_ps2_keyboard/_0365_ ), .Z(\u_ps2_keyboard/_0172_ ) );
MUX2_X1 \u_ps2_keyboard/_0654_ ( .A(\u_ps2_keyboard/_0261_ ), .B(\u_ps2_keyboard/_0200_ ), .S(\u_ps2_keyboard/_0365_ ), .Z(\u_ps2_keyboard/_0173_ ) );
NAND2_X1 \u_ps2_keyboard/_0655_ ( .A1(\u_ps2_keyboard/_0337_ ), .A2(\u_ps2_keyboard/_0361_ ), .ZN(\u_ps2_keyboard/_0366_ ) );
MUX2_X1 \u_ps2_keyboard/_0656_ ( .A(\u_ps2_keyboard/_0432_ ), .B(\u_ps2_keyboard/_0194_ ), .S(\u_ps2_keyboard/_0366_ ), .Z(\u_ps2_keyboard/_0098_ ) );
NAND2_X1 \u_ps2_keyboard/_0657_ ( .A1(\u_ps2_keyboard/_0323_ ), .A2(\u_ps2_keyboard/_0361_ ), .ZN(\u_ps2_keyboard/_0367_ ) );
MUX2_X1 \u_ps2_keyboard/_0658_ ( .A(\u_ps2_keyboard/_0432_ ), .B(\u_ps2_keyboard/_0193_ ), .S(\u_ps2_keyboard/_0367_ ), .Z(\u_ps2_keyboard/_0097_ ) );
INV_X1 \u_ps2_keyboard/_0659_ ( .A(\u_ps2_keyboard/_0184_ ), .ZN(\u_ps2_keyboard/_0368_ ) );
AND2_X1 \u_ps2_keyboard/_0660_ ( .A1(\u_ps2_keyboard/_0320_ ), .A2(\u_ps2_keyboard/_0437_ ), .ZN(\u_ps2_keyboard/_0369_ ) );
NAND3_X4 \u_ps2_keyboard/_0661_ ( .A1(\u_ps2_keyboard/_0356_ ), .A2(\u_ps2_keyboard/_0368_ ), .A3(\u_ps2_keyboard/_0369_ ), .ZN(\u_ps2_keyboard/_0370_ ) );
INV_X1 \u_ps2_keyboard/_0662_ ( .A(\u_ps2_keyboard/_0447_ ), .ZN(\u_ps2_keyboard/_0371_ ) );
NAND2_X1 \u_ps2_keyboard/_0663_ ( .A1(\u_ps2_keyboard/_0371_ ), .A2(\u_ps2_keyboard/_0448_ ), .ZN(\u_ps2_keyboard/_0372_ ) );
NOR2_X4 \u_ps2_keyboard/_0664_ ( .A1(\u_ps2_keyboard/_0370_ ), .A2(\u_ps2_keyboard/_0372_ ), .ZN(\u_ps2_keyboard/_0373_ ) );
MUX2_X1 \u_ps2_keyboard/_0665_ ( .A(\u_ps2_keyboard/_0246_ ), .B(\u_ps2_keyboard/_0193_ ), .S(\u_ps2_keyboard/_0373_ ), .Z(\u_ps2_keyboard/_0158_ ) );
MUX2_X1 \u_ps2_keyboard/_0666_ ( .A(\u_ps2_keyboard/_0247_ ), .B(\u_ps2_keyboard/_0194_ ), .S(\u_ps2_keyboard/_0373_ ), .Z(\u_ps2_keyboard/_0159_ ) );
MUX2_X1 \u_ps2_keyboard/_0667_ ( .A(\u_ps2_keyboard/_0248_ ), .B(\u_ps2_keyboard/_0195_ ), .S(\u_ps2_keyboard/_0373_ ), .Z(\u_ps2_keyboard/_0160_ ) );
MUX2_X1 \u_ps2_keyboard/_0668_ ( .A(\u_ps2_keyboard/_0249_ ), .B(\u_ps2_keyboard/_0196_ ), .S(\u_ps2_keyboard/_0373_ ), .Z(\u_ps2_keyboard/_0161_ ) );
MUX2_X1 \u_ps2_keyboard/_0669_ ( .A(\u_ps2_keyboard/_0250_ ), .B(\u_ps2_keyboard/_0197_ ), .S(\u_ps2_keyboard/_0373_ ), .Z(\u_ps2_keyboard/_0162_ ) );
MUX2_X1 \u_ps2_keyboard/_0670_ ( .A(\u_ps2_keyboard/_0251_ ), .B(\u_ps2_keyboard/_0198_ ), .S(\u_ps2_keyboard/_0373_ ), .Z(\u_ps2_keyboard/_0163_ ) );
MUX2_X1 \u_ps2_keyboard/_0671_ ( .A(\u_ps2_keyboard/_0252_ ), .B(\u_ps2_keyboard/_0199_ ), .S(\u_ps2_keyboard/_0373_ ), .Z(\u_ps2_keyboard/_0164_ ) );
MUX2_X1 \u_ps2_keyboard/_0672_ ( .A(\u_ps2_keyboard/_0253_ ), .B(\u_ps2_keyboard/_0200_ ), .S(\u_ps2_keyboard/_0373_ ), .Z(\u_ps2_keyboard/_0165_ ) );
NAND2_X1 \u_ps2_keyboard/_0673_ ( .A1(\u_ps2_keyboard/_0329_ ), .A2(\u_ps2_keyboard/_0361_ ), .ZN(\u_ps2_keyboard/_0374_ ) );
MUX2_X1 \u_ps2_keyboard/_0674_ ( .A(\u_ps2_keyboard/_0432_ ), .B(\u_ps2_keyboard/_0192_ ), .S(\u_ps2_keyboard/_0374_ ), .Z(\u_ps2_keyboard/_0096_ ) );
AND2_X4 \u_ps2_keyboard/_0675_ ( .A1(\u_ps2_keyboard/_0356_ ), .A2(\u_ps2_keyboard/_0369_ ), .ZN(\u_ps2_keyboard/_0375_ ) );
NAND2_X4 \u_ps2_keyboard/_0676_ ( .A1(\u_ps2_keyboard/_0375_ ), .A2(\u_ps2_keyboard/_0363_ ), .ZN(\u_ps2_keyboard/_0376_ ) );
NOR2_X4 \u_ps2_keyboard/_0677_ ( .A1(\u_ps2_keyboard/_0376_ ), .A2(\u_ps2_keyboard/_0372_ ), .ZN(\u_ps2_keyboard/_0377_ ) );
MUX2_X1 \u_ps2_keyboard/_0678_ ( .A(\u_ps2_keyboard/_0238_ ), .B(\u_ps2_keyboard/_0193_ ), .S(\u_ps2_keyboard/_0377_ ), .Z(\u_ps2_keyboard/_0150_ ) );
MUX2_X1 \u_ps2_keyboard/_0679_ ( .A(\u_ps2_keyboard/_0239_ ), .B(\u_ps2_keyboard/_0194_ ), .S(\u_ps2_keyboard/_0377_ ), .Z(\u_ps2_keyboard/_0151_ ) );
MUX2_X1 \u_ps2_keyboard/_0680_ ( .A(\u_ps2_keyboard/_0240_ ), .B(\u_ps2_keyboard/_0195_ ), .S(\u_ps2_keyboard/_0377_ ), .Z(\u_ps2_keyboard/_0152_ ) );
MUX2_X1 \u_ps2_keyboard/_0681_ ( .A(\u_ps2_keyboard/_0241_ ), .B(\u_ps2_keyboard/_0196_ ), .S(\u_ps2_keyboard/_0377_ ), .Z(\u_ps2_keyboard/_0153_ ) );
MUX2_X1 \u_ps2_keyboard/_0682_ ( .A(\u_ps2_keyboard/_0242_ ), .B(\u_ps2_keyboard/_0197_ ), .S(\u_ps2_keyboard/_0377_ ), .Z(\u_ps2_keyboard/_0154_ ) );
MUX2_X1 \u_ps2_keyboard/_0683_ ( .A(\u_ps2_keyboard/_0243_ ), .B(\u_ps2_keyboard/_0198_ ), .S(\u_ps2_keyboard/_0377_ ), .Z(\u_ps2_keyboard/_0155_ ) );
MUX2_X1 \u_ps2_keyboard/_0684_ ( .A(\u_ps2_keyboard/_0244_ ), .B(\u_ps2_keyboard/_0199_ ), .S(\u_ps2_keyboard/_0377_ ), .Z(\u_ps2_keyboard/_0156_ ) );
MUX2_X1 \u_ps2_keyboard/_0685_ ( .A(\u_ps2_keyboard/_0245_ ), .B(\u_ps2_keyboard/_0200_ ), .S(\u_ps2_keyboard/_0377_ ), .Z(\u_ps2_keyboard/_0157_ ) );
INV_X1 \u_ps2_keyboard/_0686_ ( .A(\u_ps2_keyboard/_0448_ ), .ZN(\u_ps2_keyboard/_0378_ ) );
NAND2_X1 \u_ps2_keyboard/_0687_ ( .A1(\u_ps2_keyboard/_0378_ ), .A2(\u_ps2_keyboard/_0447_ ), .ZN(\u_ps2_keyboard/_0379_ ) );
NOR2_X4 \u_ps2_keyboard/_0688_ ( .A1(\u_ps2_keyboard/_0370_ ), .A2(\u_ps2_keyboard/_0379_ ), .ZN(\u_ps2_keyboard/_0380_ ) );
MUX2_X1 \u_ps2_keyboard/_0689_ ( .A(\u_ps2_keyboard/_0230_ ), .B(\u_ps2_keyboard/_0193_ ), .S(\u_ps2_keyboard/_0380_ ), .Z(\u_ps2_keyboard/_0142_ ) );
MUX2_X1 \u_ps2_keyboard/_0690_ ( .A(\u_ps2_keyboard/_0231_ ), .B(\u_ps2_keyboard/_0194_ ), .S(\u_ps2_keyboard/_0380_ ), .Z(\u_ps2_keyboard/_0143_ ) );
MUX2_X1 \u_ps2_keyboard/_0691_ ( .A(\u_ps2_keyboard/_0232_ ), .B(\u_ps2_keyboard/_0195_ ), .S(\u_ps2_keyboard/_0380_ ), .Z(\u_ps2_keyboard/_0144_ ) );
MUX2_X1 \u_ps2_keyboard/_0692_ ( .A(\u_ps2_keyboard/_0233_ ), .B(\u_ps2_keyboard/_0196_ ), .S(\u_ps2_keyboard/_0380_ ), .Z(\u_ps2_keyboard/_0145_ ) );
MUX2_X1 \u_ps2_keyboard/_0693_ ( .A(\u_ps2_keyboard/_0234_ ), .B(\u_ps2_keyboard/_0197_ ), .S(\u_ps2_keyboard/_0380_ ), .Z(\u_ps2_keyboard/_0146_ ) );
MUX2_X1 \u_ps2_keyboard/_0694_ ( .A(\u_ps2_keyboard/_0235_ ), .B(\u_ps2_keyboard/_0198_ ), .S(\u_ps2_keyboard/_0380_ ), .Z(\u_ps2_keyboard/_0147_ ) );
MUX2_X1 \u_ps2_keyboard/_0695_ ( .A(\u_ps2_keyboard/_0236_ ), .B(\u_ps2_keyboard/_0199_ ), .S(\u_ps2_keyboard/_0380_ ), .Z(\u_ps2_keyboard/_0148_ ) );
MUX2_X1 \u_ps2_keyboard/_0696_ ( .A(\u_ps2_keyboard/_0237_ ), .B(\u_ps2_keyboard/_0200_ ), .S(\u_ps2_keyboard/_0380_ ), .Z(\u_ps2_keyboard/_0149_ ) );
AND2_X1 \u_ps2_keyboard/_0697_ ( .A1(\u_ps2_keyboard/_0337_ ), .A2(\u_ps2_keyboard/_0354_ ), .ZN(\u_ps2_keyboard/_0381_ ) );
AND2_X1 \u_ps2_keyboard/_0698_ ( .A1(\u_ps2_keyboard/_0352_ ), .A2(\u_ps2_keyboard/_0381_ ), .ZN(\u_ps2_keyboard/_0382_ ) );
OAI21_X1 \u_ps2_keyboard/_0699_ ( .A(\u_ps2_keyboard/_0437_ ), .B1(\u_ps2_keyboard/_0382_ ), .B2(\u_ps2_keyboard/_0368_ ), .ZN(\u_ps2_keyboard/_0383_ ) );
AOI21_X1 \u_ps2_keyboard/_0700_ ( .A(\u_ps2_keyboard/_0383_ ), .B1(\u_ps2_keyboard/_0368_ ), .B2(\u_ps2_keyboard/_0357_ ), .ZN(\u_ps2_keyboard/_0115_ ) );
INV_X1 \u_ps2_keyboard/_0701_ ( .A(\u_ps2_keyboard/_0437_ ), .ZN(\u_ps2_keyboard/_0384_ ) );
INV_X1 \u_ps2_keyboard/_0702_ ( .A(\u_ps2_keyboard/_0356_ ), .ZN(\u_ps2_keyboard/_0385_ ) );
XNOR2_X1 \u_ps2_keyboard/_0703_ ( .A(\u_ps2_keyboard/_0447_ ), .B(\u_ps2_keyboard/_0446_ ), .ZN(\u_ps2_keyboard/_0386_ ) );
NOR2_X1 \u_ps2_keyboard/_0704_ ( .A1(\u_ps2_keyboard/_0385_ ), .A2(\u_ps2_keyboard/_0386_ ), .ZN(\u_ps2_keyboard/_0387_ ) );
INV_X1 \u_ps2_keyboard/_0705_ ( .A(\u_ps2_keyboard/_0320_ ), .ZN(\u_ps2_keyboard/_0388_ ) );
AOI21_X1 \u_ps2_keyboard/_0706_ ( .A(\u_ps2_keyboard/_0185_ ), .B1(\u_ps2_keyboard/_0352_ ), .B2(\u_ps2_keyboard/_0355_ ), .ZN(\u_ps2_keyboard/_0389_ ) );
NOR3_X1 \u_ps2_keyboard/_0707_ ( .A1(\u_ps2_keyboard/_0387_ ), .A2(\u_ps2_keyboard/_0388_ ), .A3(\u_ps2_keyboard/_0389_ ), .ZN(\u_ps2_keyboard/_0390_ ) );
AOI211_X2 \u_ps2_keyboard/_0708_ ( .A(\u_ps2_keyboard/_0384_ ), .B(\u_ps2_keyboard/_0390_ ), .C1(\u_ps2_keyboard/_0185_ ), .C2(\u_ps2_keyboard/_0388_ ), .ZN(\u_ps2_keyboard/_0116_ ) );
NAND2_X1 \u_ps2_keyboard/_0709_ ( .A1(\u_ps2_keyboard/_0447_ ), .A2(\u_ps2_keyboard/_0446_ ), .ZN(\u_ps2_keyboard/_0391_ ) );
XNOR2_X1 \u_ps2_keyboard/_0710_ ( .A(\u_ps2_keyboard/_0391_ ), .B(\u_ps2_keyboard/_0186_ ), .ZN(\u_ps2_keyboard/_0392_ ) );
AND4_X1 \u_ps2_keyboard/_0711_ ( .A1(\u_ps2_keyboard/_0351_ ), .A2(\u_ps2_keyboard/_0350_ ), .A3(\u_ps2_keyboard/_0381_ ), .A4(\u_ps2_keyboard/_0392_ ), .ZN(\u_ps2_keyboard/_0393_ ) );
INV_X1 \u_ps2_keyboard/_0712_ ( .A(\u_ps2_keyboard/_0382_ ), .ZN(\u_ps2_keyboard/_0394_ ) );
AOI211_X4 \u_ps2_keyboard/_0713_ ( .A(\u_ps2_keyboard/_0384_ ), .B(\u_ps2_keyboard/_0393_ ), .C1(\u_ps2_keyboard/_0394_ ), .C2(\u_ps2_keyboard/_0186_ ), .ZN(\u_ps2_keyboard/_0117_ ) );
XNOR2_X1 \u_ps2_keyboard/_0714_ ( .A(\u_ps2_keyboard/_0433_ ), .B(\u_ps2_keyboard/_0428_ ), .ZN(\u_ps2_keyboard/_0395_ ) );
NAND2_X1 \u_ps2_keyboard/_0715_ ( .A1(\u_ps2_keyboard/_0395_ ), .A2(\u_ps2_keyboard/_0436_ ), .ZN(\u_ps2_keyboard/_0396_ ) );
OR2_X1 \u_ps2_keyboard/_0716_ ( .A1(\u_ps2_keyboard/_0187_ ), .A2(\u_ps2_keyboard/_0436_ ), .ZN(\u_ps2_keyboard/_0397_ ) );
AOI21_X1 \u_ps2_keyboard/_0717_ ( .A(\u_ps2_keyboard/_0384_ ), .B1(\u_ps2_keyboard/_0396_ ), .B2(\u_ps2_keyboard/_0397_ ), .ZN(\u_ps2_keyboard/_0111_ ) );
XOR2_X1 \u_ps2_keyboard/_0718_ ( .A(\u_ps2_keyboard/_0433_ ), .B(\u_ps2_keyboard/_0434_ ), .Z(\u_ps2_keyboard/_0398_ ) );
INV_X1 \u_ps2_keyboard/_0719_ ( .A(\u_ps2_keyboard/_0428_ ), .ZN(\u_ps2_keyboard/_0399_ ) );
NAND2_X1 \u_ps2_keyboard/_0720_ ( .A1(\u_ps2_keyboard/_0399_ ), .A2(\u_ps2_keyboard/_0436_ ), .ZN(\u_ps2_keyboard/_0400_ ) );
NOR2_X1 \u_ps2_keyboard/_0721_ ( .A1(\u_ps2_keyboard/_0398_ ), .A2(\u_ps2_keyboard/_0400_ ), .ZN(\u_ps2_keyboard/_0401_ ) );
AOI211_X4 \u_ps2_keyboard/_0722_ ( .A(\u_ps2_keyboard/_0384_ ), .B(\u_ps2_keyboard/_0401_ ), .C1(\u_ps2_keyboard/_0183_ ), .C2(\u_ps2_keyboard/_0400_ ), .ZN(\u_ps2_keyboard/_0112_ ) );
NAND2_X1 \u_ps2_keyboard/_0723_ ( .A1(\u_ps2_keyboard/_0433_ ), .A2(\u_ps2_keyboard/_0434_ ), .ZN(\u_ps2_keyboard/_0402_ ) );
XNOR2_X1 \u_ps2_keyboard/_0724_ ( .A(\u_ps2_keyboard/_0402_ ), .B(\u_ps2_keyboard/_0182_ ), .ZN(\u_ps2_keyboard/_0403_ ) );
AND3_X1 \u_ps2_keyboard/_0725_ ( .A1(\u_ps2_keyboard/_0403_ ), .A2(\u_ps2_keyboard/_0399_ ), .A3(\u_ps2_keyboard/_0436_ ), .ZN(\u_ps2_keyboard/_0404_ ) );
AOI211_X4 \u_ps2_keyboard/_0726_ ( .A(\u_ps2_keyboard/_0384_ ), .B(\u_ps2_keyboard/_0404_ ), .C1(\u_ps2_keyboard/_0182_ ), .C2(\u_ps2_keyboard/_0400_ ), .ZN(\u_ps2_keyboard/_0113_ ) );
NOR2_X4 \u_ps2_keyboard/_0727_ ( .A1(\u_ps2_keyboard/_0376_ ), .A2(\u_ps2_keyboard/_0379_ ), .ZN(\u_ps2_keyboard/_0405_ ) );
MUX2_X1 \u_ps2_keyboard/_0728_ ( .A(\u_ps2_keyboard/_0222_ ), .B(\u_ps2_keyboard/_0193_ ), .S(\u_ps2_keyboard/_0405_ ), .Z(\u_ps2_keyboard/_0134_ ) );
MUX2_X1 \u_ps2_keyboard/_0729_ ( .A(\u_ps2_keyboard/_0223_ ), .B(\u_ps2_keyboard/_0194_ ), .S(\u_ps2_keyboard/_0405_ ), .Z(\u_ps2_keyboard/_0135_ ) );
MUX2_X1 \u_ps2_keyboard/_0730_ ( .A(\u_ps2_keyboard/_0224_ ), .B(\u_ps2_keyboard/_0195_ ), .S(\u_ps2_keyboard/_0405_ ), .Z(\u_ps2_keyboard/_0136_ ) );
MUX2_X1 \u_ps2_keyboard/_0731_ ( .A(\u_ps2_keyboard/_0225_ ), .B(\u_ps2_keyboard/_0196_ ), .S(\u_ps2_keyboard/_0405_ ), .Z(\u_ps2_keyboard/_0137_ ) );
MUX2_X1 \u_ps2_keyboard/_0732_ ( .A(\u_ps2_keyboard/_0226_ ), .B(\u_ps2_keyboard/_0197_ ), .S(\u_ps2_keyboard/_0405_ ), .Z(\u_ps2_keyboard/_0138_ ) );
MUX2_X1 \u_ps2_keyboard/_0733_ ( .A(\u_ps2_keyboard/_0227_ ), .B(\u_ps2_keyboard/_0198_ ), .S(\u_ps2_keyboard/_0405_ ), .Z(\u_ps2_keyboard/_0139_ ) );
MUX2_X1 \u_ps2_keyboard/_0734_ ( .A(\u_ps2_keyboard/_0228_ ), .B(\u_ps2_keyboard/_0199_ ), .S(\u_ps2_keyboard/_0405_ ), .Z(\u_ps2_keyboard/_0140_ ) );
MUX2_X1 \u_ps2_keyboard/_0735_ ( .A(\u_ps2_keyboard/_0229_ ), .B(\u_ps2_keyboard/_0200_ ), .S(\u_ps2_keyboard/_0405_ ), .Z(\u_ps2_keyboard/_0141_ ) );
XNOR2_X1 \u_ps2_keyboard/_0736_ ( .A(\u_ps2_keyboard/_0320_ ), .B(\u_ps2_keyboard/_0202_ ), .ZN(\u_ps2_keyboard/_0406_ ) );
NOR3_X1 \u_ps2_keyboard/_0737_ ( .A1(\u_ps2_keyboard/_0381_ ), .A2(\u_ps2_keyboard/_0384_ ), .A3(\u_ps2_keyboard/_0406_ ), .ZN(\u_ps2_keyboard/_0106_ ) );
NOR3_X1 \u_ps2_keyboard/_0738_ ( .A1(\u_ps2_keyboard/_0322_ ), .A2(\u_ps2_keyboard/_0430_ ), .A3(\u_ps2_keyboard/_0319_ ), .ZN(\u_ps2_keyboard/_0407_ ) );
OAI211_X2 \u_ps2_keyboard/_0739_ ( .A(\u_ps2_keyboard/_0321_ ), .B(\u_ps2_keyboard/_0203_ ), .C1(\u_ps2_keyboard/_0334_ ), .C2(\u_ps2_keyboard/_0204_ ), .ZN(\u_ps2_keyboard/_0408_ ) );
AOI221_X4 \u_ps2_keyboard/_0740_ ( .A(\u_ps2_keyboard/_0384_ ), .B1(\u_ps2_keyboard/_0388_ ), .B2(\u_ps2_keyboard/_0188_ ), .C1(\u_ps2_keyboard/_0407_ ), .C2(\u_ps2_keyboard/_0408_ ), .ZN(\u_ps2_keyboard/_0107_ ) );
AND2_X1 \u_ps2_keyboard/_0741_ ( .A1(\u_ps2_keyboard/_0320_ ), .A2(\u_ps2_keyboard/_0332_ ), .ZN(\u_ps2_keyboard/_0409_ ) );
XNOR2_X1 \u_ps2_keyboard/_0742_ ( .A(\u_ps2_keyboard/_0409_ ), .B(\u_ps2_keyboard/_0189_ ), .ZN(\u_ps2_keyboard/_0410_ ) );
INV_X1 \u_ps2_keyboard/_0743_ ( .A(\u_ps2_keyboard/_0381_ ), .ZN(\u_ps2_keyboard/_0411_ ) );
AND3_X1 \u_ps2_keyboard/_0744_ ( .A1(\u_ps2_keyboard/_0410_ ), .A2(\u_ps2_keyboard/_0411_ ), .A3(\u_ps2_keyboard/_0437_ ), .ZN(\u_ps2_keyboard/_0108_ ) );
AOI221_X4 \u_ps2_keyboard/_0745_ ( .A(\u_ps2_keyboard/_0384_ ), .B1(\u_ps2_keyboard/_0333_ ), .B2(\u_ps2_keyboard/_0190_ ), .C1(\u_ps2_keyboard/_0354_ ), .C2(\u_ps2_keyboard/_0337_ ), .ZN(\u_ps2_keyboard/_0412_ ) );
OR2_X1 \u_ps2_keyboard/_0746_ ( .A1(\u_ps2_keyboard/_0333_ ), .A2(\u_ps2_keyboard/_0190_ ), .ZN(\u_ps2_keyboard/_0413_ ) );
AND2_X1 \u_ps2_keyboard/_0747_ ( .A1(\u_ps2_keyboard/_0412_ ), .A2(\u_ps2_keyboard/_0413_ ), .ZN(\u_ps2_keyboard/_0109_ ) );
NAND2_X1 \u_ps2_keyboard/_0748_ ( .A1(\u_ps2_keyboard/_0378_ ), .A2(\u_ps2_keyboard/_0371_ ), .ZN(\u_ps2_keyboard/_0414_ ) );
NOR2_X4 \u_ps2_keyboard/_0749_ ( .A1(\u_ps2_keyboard/_0370_ ), .A2(\u_ps2_keyboard/_0414_ ), .ZN(\u_ps2_keyboard/_0415_ ) );
MUX2_X1 \u_ps2_keyboard/_0750_ ( .A(\u_ps2_keyboard/_0214_ ), .B(\u_ps2_keyboard/_0193_ ), .S(\u_ps2_keyboard/_0415_ ), .Z(\u_ps2_keyboard/_0126_ ) );
MUX2_X1 \u_ps2_keyboard/_0751_ ( .A(\u_ps2_keyboard/_0215_ ), .B(\u_ps2_keyboard/_0194_ ), .S(\u_ps2_keyboard/_0415_ ), .Z(\u_ps2_keyboard/_0127_ ) );
MUX2_X1 \u_ps2_keyboard/_0752_ ( .A(\u_ps2_keyboard/_0216_ ), .B(\u_ps2_keyboard/_0195_ ), .S(\u_ps2_keyboard/_0415_ ), .Z(\u_ps2_keyboard/_0128_ ) );
MUX2_X1 \u_ps2_keyboard/_0753_ ( .A(\u_ps2_keyboard/_0217_ ), .B(\u_ps2_keyboard/_0196_ ), .S(\u_ps2_keyboard/_0415_ ), .Z(\u_ps2_keyboard/_0129_ ) );
MUX2_X1 \u_ps2_keyboard/_0754_ ( .A(\u_ps2_keyboard/_0218_ ), .B(\u_ps2_keyboard/_0197_ ), .S(\u_ps2_keyboard/_0415_ ), .Z(\u_ps2_keyboard/_0130_ ) );
MUX2_X1 \u_ps2_keyboard/_0755_ ( .A(\u_ps2_keyboard/_0219_ ), .B(\u_ps2_keyboard/_0198_ ), .S(\u_ps2_keyboard/_0415_ ), .Z(\u_ps2_keyboard/_0131_ ) );
MUX2_X1 \u_ps2_keyboard/_0756_ ( .A(\u_ps2_keyboard/_0220_ ), .B(\u_ps2_keyboard/_0199_ ), .S(\u_ps2_keyboard/_0415_ ), .Z(\u_ps2_keyboard/_0132_ ) );
MUX2_X1 \u_ps2_keyboard/_0757_ ( .A(\u_ps2_keyboard/_0221_ ), .B(\u_ps2_keyboard/_0200_ ), .S(\u_ps2_keyboard/_0415_ ), .Z(\u_ps2_keyboard/_0133_ ) );
NOR2_X4 \u_ps2_keyboard/_0758_ ( .A1(\u_ps2_keyboard/_0376_ ), .A2(\u_ps2_keyboard/_0414_ ), .ZN(\u_ps2_keyboard/_0416_ ) );
MUX2_X1 \u_ps2_keyboard/_0759_ ( .A(\u_ps2_keyboard/_0206_ ), .B(\u_ps2_keyboard/_0193_ ), .S(\u_ps2_keyboard/_0416_ ), .Z(\u_ps2_keyboard/_0118_ ) );
MUX2_X1 \u_ps2_keyboard/_0760_ ( .A(\u_ps2_keyboard/_0207_ ), .B(\u_ps2_keyboard/_0194_ ), .S(\u_ps2_keyboard/_0416_ ), .Z(\u_ps2_keyboard/_0119_ ) );
MUX2_X1 \u_ps2_keyboard/_0761_ ( .A(\u_ps2_keyboard/_0208_ ), .B(\u_ps2_keyboard/_0195_ ), .S(\u_ps2_keyboard/_0416_ ), .Z(\u_ps2_keyboard/_0120_ ) );
MUX2_X1 \u_ps2_keyboard/_0762_ ( .A(\u_ps2_keyboard/_0209_ ), .B(\u_ps2_keyboard/_0196_ ), .S(\u_ps2_keyboard/_0416_ ), .Z(\u_ps2_keyboard/_0121_ ) );
MUX2_X1 \u_ps2_keyboard/_0763_ ( .A(\u_ps2_keyboard/_0210_ ), .B(\u_ps2_keyboard/_0197_ ), .S(\u_ps2_keyboard/_0416_ ), .Z(\u_ps2_keyboard/_0122_ ) );
MUX2_X1 \u_ps2_keyboard/_0764_ ( .A(\u_ps2_keyboard/_0211_ ), .B(\u_ps2_keyboard/_0198_ ), .S(\u_ps2_keyboard/_0416_ ), .Z(\u_ps2_keyboard/_0123_ ) );
MUX2_X1 \u_ps2_keyboard/_0765_ ( .A(\u_ps2_keyboard/_0212_ ), .B(\u_ps2_keyboard/_0199_ ), .S(\u_ps2_keyboard/_0416_ ), .Z(\u_ps2_keyboard/_0124_ ) );
MUX2_X1 \u_ps2_keyboard/_0766_ ( .A(\u_ps2_keyboard/_0213_ ), .B(\u_ps2_keyboard/_0200_ ), .S(\u_ps2_keyboard/_0416_ ), .Z(\u_ps2_keyboard/_0125_ ) );
XNOR2_X1 \u_ps2_keyboard/_0767_ ( .A(\u_ps2_keyboard/_0398_ ), .B(\u_ps2_keyboard/_0185_ ), .ZN(\u_ps2_keyboard/_0417_ ) );
XNOR2_X1 \u_ps2_keyboard/_0768_ ( .A(\u_ps2_keyboard/_0433_ ), .B(\u_ps2_keyboard/_0446_ ), .ZN(\u_ps2_keyboard/_0418_ ) );
NOR3_X1 \u_ps2_keyboard/_0769_ ( .A1(\u_ps2_keyboard/_0417_ ), .A2(\u_ps2_keyboard/_0428_ ), .A3(\u_ps2_keyboard/_0418_ ), .ZN(\u_ps2_keyboard/_0419_ ) );
XNOR2_X1 \u_ps2_keyboard/_0770_ ( .A(\u_ps2_keyboard/_0403_ ), .B(\u_ps2_keyboard/_0186_ ), .ZN(\u_ps2_keyboard/_0420_ ) );
NAND2_X1 \u_ps2_keyboard/_0771_ ( .A1(\u_ps2_keyboard/_0419_ ), .A2(\u_ps2_keyboard/_0420_ ), .ZN(\u_ps2_keyboard/_0421_ ) );
AND3_X1 \u_ps2_keyboard/_0772_ ( .A1(\u_ps2_keyboard/_0421_ ), .A2(\u_ps2_keyboard/_0437_ ), .A3(\u_ps2_keyboard/_0436_ ), .ZN(\u_ps2_keyboard/_0422_ ) );
OR2_X1 \u_ps2_keyboard/_0773_ ( .A1(\u_ps2_keyboard/_0375_ ), .A2(\u_ps2_keyboard/_0422_ ), .ZN(\u_ps2_keyboard/_0114_ ) );
XOR2_X1 \u_ps2_keyboard/_0774_ ( .A(\u_ps2_keyboard/_0392_ ), .B(\u_ps2_keyboard/_0182_ ), .Z(\u_ps2_keyboard/_0423_ ) );
XOR2_X1 \u_ps2_keyboard/_0775_ ( .A(\u_ps2_keyboard/_0386_ ), .B(\u_ps2_keyboard/_0183_ ), .Z(\u_ps2_keyboard/_0424_ ) );
NOR3_X1 \u_ps2_keyboard/_0776_ ( .A1(\u_ps2_keyboard/_0423_ ), .A2(\u_ps2_keyboard/_0418_ ), .A3(\u_ps2_keyboard/_0424_ ), .ZN(\u_ps2_keyboard/_0425_ ) );
NAND3_X1 \u_ps2_keyboard/_0777_ ( .A1(\u_ps2_keyboard/_0350_ ), .A2(\u_ps2_keyboard/_0351_ ), .A3(\u_ps2_keyboard/_0425_ ), .ZN(\u_ps2_keyboard/_0426_ ) );
NOR2_X1 \u_ps2_keyboard/_0778_ ( .A1(\u_ps2_keyboard/_0411_ ), .A2(\u_ps2_keyboard/_0429_ ), .ZN(\u_ps2_keyboard/_0427_ ) );
AOI221_X4 \u_ps2_keyboard/_0779_ ( .A(\u_ps2_keyboard/_0384_ ), .B1(\u_ps2_keyboard/_0191_ ), .B2(\u_ps2_keyboard/_0411_ ), .C1(\u_ps2_keyboard/_0426_ ), .C2(\u_ps2_keyboard/_0427_ ), .ZN(\u_ps2_keyboard/_0110_ ) );
BUF_X1 \u_ps2_keyboard/_0780_ ( .A(\u_ps2_keyboard/fifo[0][0] ), .Z(\u_ps2_keyboard/_0206_ ) );
BUF_X1 \u_ps2_keyboard/_0781_ ( .A(\u_ps2_keyboard/fifo[1][0] ), .Z(\u_ps2_keyboard/_0214_ ) );
BUF_X1 \u_ps2_keyboard/_0782_ ( .A(\u_ps2_keyboard/r_ptr [0] ), .Z(\u_ps2_keyboard/_0433_ ) );
BUF_X1 \u_ps2_keyboard/_0783_ ( .A(\u_ps2_keyboard/fifo[2][0] ), .Z(\u_ps2_keyboard/_0222_ ) );
BUF_X1 \u_ps2_keyboard/_0784_ ( .A(\u_ps2_keyboard/fifo[3][0] ), .Z(\u_ps2_keyboard/_0230_ ) );
BUF_X1 \u_ps2_keyboard/_0785_ ( .A(\u_ps2_keyboard/r_ptr [1] ), .Z(\u_ps2_keyboard/_0434_ ) );
BUF_X1 \u_ps2_keyboard/_0786_ ( .A(\u_ps2_keyboard/fifo[4][0] ), .Z(\u_ps2_keyboard/_0238_ ) );
BUF_X1 \u_ps2_keyboard/_0787_ ( .A(\u_ps2_keyboard/fifo[5][0] ), .Z(\u_ps2_keyboard/_0246_ ) );
BUF_X1 \u_ps2_keyboard/_0788_ ( .A(\u_ps2_keyboard/fifo[6][0] ), .Z(\u_ps2_keyboard/_0254_ ) );
BUF_X1 \u_ps2_keyboard/_0789_ ( .A(\u_ps2_keyboard/fifo[7][0] ), .Z(\u_ps2_keyboard/_0262_ ) );
BUF_X1 \u_ps2_keyboard/_0790_ ( .A(\u_ps2_keyboard/r_ptr [2] ), .Z(\u_ps2_keyboard/_0435_ ) );
BUF_X1 \u_ps2_keyboard/_0791_ ( .A(\u_ps2_keyboard/_0438_ ), .Z(\scan_code [0] ) );
BUF_X1 \u_ps2_keyboard/_0792_ ( .A(\u_ps2_keyboard/fifo[0][1] ), .Z(\u_ps2_keyboard/_0207_ ) );
BUF_X1 \u_ps2_keyboard/_0793_ ( .A(\u_ps2_keyboard/fifo[1][1] ), .Z(\u_ps2_keyboard/_0215_ ) );
BUF_X1 \u_ps2_keyboard/_0794_ ( .A(\u_ps2_keyboard/fifo[2][1] ), .Z(\u_ps2_keyboard/_0223_ ) );
BUF_X1 \u_ps2_keyboard/_0795_ ( .A(\u_ps2_keyboard/fifo[3][1] ), .Z(\u_ps2_keyboard/_0231_ ) );
BUF_X1 \u_ps2_keyboard/_0796_ ( .A(\u_ps2_keyboard/fifo[4][1] ), .Z(\u_ps2_keyboard/_0239_ ) );
BUF_X1 \u_ps2_keyboard/_0797_ ( .A(\u_ps2_keyboard/fifo[5][1] ), .Z(\u_ps2_keyboard/_0247_ ) );
BUF_X1 \u_ps2_keyboard/_0798_ ( .A(\u_ps2_keyboard/fifo[6][1] ), .Z(\u_ps2_keyboard/_0255_ ) );
BUF_X1 \u_ps2_keyboard/_0799_ ( .A(\u_ps2_keyboard/fifo[7][1] ), .Z(\u_ps2_keyboard/_0263_ ) );
BUF_X1 \u_ps2_keyboard/_0800_ ( .A(\u_ps2_keyboard/_0439_ ), .Z(\scan_code [1] ) );
BUF_X1 \u_ps2_keyboard/_0801_ ( .A(\u_ps2_keyboard/fifo[0][2] ), .Z(\u_ps2_keyboard/_0208_ ) );
BUF_X1 \u_ps2_keyboard/_0802_ ( .A(\u_ps2_keyboard/fifo[1][2] ), .Z(\u_ps2_keyboard/_0216_ ) );
BUF_X1 \u_ps2_keyboard/_0803_ ( .A(\u_ps2_keyboard/fifo[2][2] ), .Z(\u_ps2_keyboard/_0224_ ) );
BUF_X1 \u_ps2_keyboard/_0804_ ( .A(\u_ps2_keyboard/fifo[3][2] ), .Z(\u_ps2_keyboard/_0232_ ) );
BUF_X1 \u_ps2_keyboard/_0805_ ( .A(\u_ps2_keyboard/fifo[4][2] ), .Z(\u_ps2_keyboard/_0240_ ) );
BUF_X1 \u_ps2_keyboard/_0806_ ( .A(\u_ps2_keyboard/fifo[5][2] ), .Z(\u_ps2_keyboard/_0248_ ) );
BUF_X1 \u_ps2_keyboard/_0807_ ( .A(\u_ps2_keyboard/fifo[6][2] ), .Z(\u_ps2_keyboard/_0256_ ) );
BUF_X1 \u_ps2_keyboard/_0808_ ( .A(\u_ps2_keyboard/fifo[7][2] ), .Z(\u_ps2_keyboard/_0264_ ) );
BUF_X1 \u_ps2_keyboard/_0809_ ( .A(\u_ps2_keyboard/_0440_ ), .Z(\scan_code [2] ) );
BUF_X1 \u_ps2_keyboard/_0810_ ( .A(\u_ps2_keyboard/fifo[0][3] ), .Z(\u_ps2_keyboard/_0209_ ) );
BUF_X1 \u_ps2_keyboard/_0811_ ( .A(\u_ps2_keyboard/fifo[1][3] ), .Z(\u_ps2_keyboard/_0217_ ) );
BUF_X1 \u_ps2_keyboard/_0812_ ( .A(\u_ps2_keyboard/fifo[2][3] ), .Z(\u_ps2_keyboard/_0225_ ) );
BUF_X1 \u_ps2_keyboard/_0813_ ( .A(\u_ps2_keyboard/fifo[3][3] ), .Z(\u_ps2_keyboard/_0233_ ) );
BUF_X1 \u_ps2_keyboard/_0814_ ( .A(\u_ps2_keyboard/fifo[4][3] ), .Z(\u_ps2_keyboard/_0241_ ) );
BUF_X1 \u_ps2_keyboard/_0815_ ( .A(\u_ps2_keyboard/fifo[5][3] ), .Z(\u_ps2_keyboard/_0249_ ) );
BUF_X1 \u_ps2_keyboard/_0816_ ( .A(\u_ps2_keyboard/fifo[6][3] ), .Z(\u_ps2_keyboard/_0257_ ) );
BUF_X1 \u_ps2_keyboard/_0817_ ( .A(\u_ps2_keyboard/fifo[7][3] ), .Z(\u_ps2_keyboard/_0265_ ) );
BUF_X1 \u_ps2_keyboard/_0818_ ( .A(\u_ps2_keyboard/_0441_ ), .Z(\scan_code [3] ) );
BUF_X1 \u_ps2_keyboard/_0819_ ( .A(\u_ps2_keyboard/fifo[0][4] ), .Z(\u_ps2_keyboard/_0210_ ) );
BUF_X1 \u_ps2_keyboard/_0820_ ( .A(\u_ps2_keyboard/fifo[1][4] ), .Z(\u_ps2_keyboard/_0218_ ) );
BUF_X1 \u_ps2_keyboard/_0821_ ( .A(\u_ps2_keyboard/fifo[2][4] ), .Z(\u_ps2_keyboard/_0226_ ) );
BUF_X1 \u_ps2_keyboard/_0822_ ( .A(\u_ps2_keyboard/fifo[3][4] ), .Z(\u_ps2_keyboard/_0234_ ) );
BUF_X1 \u_ps2_keyboard/_0823_ ( .A(\u_ps2_keyboard/fifo[4][4] ), .Z(\u_ps2_keyboard/_0242_ ) );
BUF_X1 \u_ps2_keyboard/_0824_ ( .A(\u_ps2_keyboard/fifo[5][4] ), .Z(\u_ps2_keyboard/_0250_ ) );
BUF_X1 \u_ps2_keyboard/_0825_ ( .A(\u_ps2_keyboard/fifo[6][4] ), .Z(\u_ps2_keyboard/_0258_ ) );
BUF_X1 \u_ps2_keyboard/_0826_ ( .A(\u_ps2_keyboard/fifo[7][4] ), .Z(\u_ps2_keyboard/_0266_ ) );
BUF_X1 \u_ps2_keyboard/_0827_ ( .A(\u_ps2_keyboard/_0442_ ), .Z(\scan_code [4] ) );
BUF_X1 \u_ps2_keyboard/_0828_ ( .A(\u_ps2_keyboard/fifo[0][5] ), .Z(\u_ps2_keyboard/_0211_ ) );
BUF_X1 \u_ps2_keyboard/_0829_ ( .A(\u_ps2_keyboard/fifo[1][5] ), .Z(\u_ps2_keyboard/_0219_ ) );
BUF_X1 \u_ps2_keyboard/_0830_ ( .A(\u_ps2_keyboard/fifo[2][5] ), .Z(\u_ps2_keyboard/_0227_ ) );
BUF_X1 \u_ps2_keyboard/_0831_ ( .A(\u_ps2_keyboard/fifo[3][5] ), .Z(\u_ps2_keyboard/_0235_ ) );
BUF_X1 \u_ps2_keyboard/_0832_ ( .A(\u_ps2_keyboard/fifo[4][5] ), .Z(\u_ps2_keyboard/_0243_ ) );
BUF_X1 \u_ps2_keyboard/_0833_ ( .A(\u_ps2_keyboard/fifo[5][5] ), .Z(\u_ps2_keyboard/_0251_ ) );
BUF_X1 \u_ps2_keyboard/_0834_ ( .A(\u_ps2_keyboard/fifo[6][5] ), .Z(\u_ps2_keyboard/_0259_ ) );
BUF_X1 \u_ps2_keyboard/_0835_ ( .A(\u_ps2_keyboard/fifo[7][5] ), .Z(\u_ps2_keyboard/_0267_ ) );
BUF_X1 \u_ps2_keyboard/_0836_ ( .A(\u_ps2_keyboard/_0443_ ), .Z(\scan_code [5] ) );
BUF_X1 \u_ps2_keyboard/_0837_ ( .A(\u_ps2_keyboard/fifo[0][6] ), .Z(\u_ps2_keyboard/_0212_ ) );
BUF_X1 \u_ps2_keyboard/_0838_ ( .A(\u_ps2_keyboard/fifo[1][6] ), .Z(\u_ps2_keyboard/_0220_ ) );
BUF_X1 \u_ps2_keyboard/_0839_ ( .A(\u_ps2_keyboard/fifo[2][6] ), .Z(\u_ps2_keyboard/_0228_ ) );
BUF_X1 \u_ps2_keyboard/_0840_ ( .A(\u_ps2_keyboard/fifo[3][6] ), .Z(\u_ps2_keyboard/_0236_ ) );
BUF_X1 \u_ps2_keyboard/_0841_ ( .A(\u_ps2_keyboard/fifo[4][6] ), .Z(\u_ps2_keyboard/_0244_ ) );
BUF_X1 \u_ps2_keyboard/_0842_ ( .A(\u_ps2_keyboard/fifo[5][6] ), .Z(\u_ps2_keyboard/_0252_ ) );
BUF_X1 \u_ps2_keyboard/_0843_ ( .A(\u_ps2_keyboard/fifo[6][6] ), .Z(\u_ps2_keyboard/_0260_ ) );
BUF_X1 \u_ps2_keyboard/_0844_ ( .A(\u_ps2_keyboard/fifo[7][6] ), .Z(\u_ps2_keyboard/_0268_ ) );
BUF_X1 \u_ps2_keyboard/_0845_ ( .A(\u_ps2_keyboard/_0444_ ), .Z(\scan_code [6] ) );
BUF_X1 \u_ps2_keyboard/_0846_ ( .A(\u_ps2_keyboard/fifo[0][7] ), .Z(\u_ps2_keyboard/_0213_ ) );
BUF_X1 \u_ps2_keyboard/_0847_ ( .A(\u_ps2_keyboard/fifo[1][7] ), .Z(\u_ps2_keyboard/_0221_ ) );
BUF_X1 \u_ps2_keyboard/_0848_ ( .A(\u_ps2_keyboard/fifo[2][7] ), .Z(\u_ps2_keyboard/_0229_ ) );
BUF_X1 \u_ps2_keyboard/_0849_ ( .A(\u_ps2_keyboard/fifo[3][7] ), .Z(\u_ps2_keyboard/_0237_ ) );
BUF_X1 \u_ps2_keyboard/_0850_ ( .A(\u_ps2_keyboard/fifo[4][7] ), .Z(\u_ps2_keyboard/_0245_ ) );
BUF_X1 \u_ps2_keyboard/_0851_ ( .A(\u_ps2_keyboard/fifo[5][7] ), .Z(\u_ps2_keyboard/_0253_ ) );
BUF_X1 \u_ps2_keyboard/_0852_ ( .A(\u_ps2_keyboard/fifo[6][7] ), .Z(\u_ps2_keyboard/_0261_ ) );
BUF_X1 \u_ps2_keyboard/_0853_ ( .A(\u_ps2_keyboard/fifo[7][7] ), .Z(\u_ps2_keyboard/_0269_ ) );
BUF_X1 \u_ps2_keyboard/_0854_ ( .A(\u_ps2_keyboard/_0445_ ), .Z(\scan_code [7] ) );
BUF_X1 \u_ps2_keyboard/_0855_ ( .A(rst_n ), .Z(\u_ps2_keyboard/_0437_ ) );
BUF_X1 \u_ps2_keyboard/_0856_ ( .A(\u_ps2_keyboard/ps2_clk_sync [1] ), .Z(\u_ps2_keyboard/_0430_ ) );
BUF_X1 \u_ps2_keyboard/_0857_ ( .A(\u_ps2_keyboard/ps2_clk_sync [2] ), .Z(\u_ps2_keyboard/_0431_ ) );
BUF_X1 \u_ps2_keyboard/_0858_ ( .A(\u_ps2_keyboard/count [2] ), .Z(\u_ps2_keyboard/_0204_ ) );
BUF_X1 \u_ps2_keyboard/_0859_ ( .A(\u_ps2_keyboard/count [3] ), .Z(\u_ps2_keyboard/_0205_ ) );
BUF_X1 \u_ps2_keyboard/_0860_ ( .A(\u_ps2_keyboard/count [0] ), .Z(\u_ps2_keyboard/_0202_ ) );
BUF_X1 \u_ps2_keyboard/_0861_ ( .A(\u_ps2_keyboard/count [1] ), .Z(\u_ps2_keyboard/_0203_ ) );
BUF_X1 \u_ps2_keyboard/_0862_ ( .A(ps2_data ), .Z(\u_ps2_keyboard/_0432_ ) );
BUF_X1 \u_ps2_keyboard/_0863_ ( .A(\u_ps2_keyboard/buffer [9] ), .Z(\u_ps2_keyboard/_0201_ ) );
BUF_X1 \u_ps2_keyboard/_0864_ ( .A(\u_ps2_keyboard/_0105_ ), .Z(\u_ps2_keyboard/_0009_ ) );
BUF_X1 \u_ps2_keyboard/_0865_ ( .A(\u_ps2_keyboard/buffer [8] ), .Z(\u_ps2_keyboard/_0200_ ) );
BUF_X1 \u_ps2_keyboard/_0866_ ( .A(\u_ps2_keyboard/_0104_ ), .Z(\u_ps2_keyboard/_0008_ ) );
BUF_X1 \u_ps2_keyboard/_0867_ ( .A(\u_ps2_keyboard/buffer [7] ), .Z(\u_ps2_keyboard/_0199_ ) );
BUF_X1 \u_ps2_keyboard/_0868_ ( .A(\u_ps2_keyboard/_0103_ ), .Z(\u_ps2_keyboard/_0007_ ) );
BUF_X1 \u_ps2_keyboard/_0869_ ( .A(\u_ps2_keyboard/buffer [6] ), .Z(\u_ps2_keyboard/_0198_ ) );
BUF_X1 \u_ps2_keyboard/_0870_ ( .A(\u_ps2_keyboard/_0102_ ), .Z(\u_ps2_keyboard/_0006_ ) );
BUF_X1 \u_ps2_keyboard/_0871_ ( .A(\u_ps2_keyboard/buffer [5] ), .Z(\u_ps2_keyboard/_0197_ ) );
BUF_X1 \u_ps2_keyboard/_0872_ ( .A(\u_ps2_keyboard/_0101_ ), .Z(\u_ps2_keyboard/_0005_ ) );
BUF_X1 \u_ps2_keyboard/_0873_ ( .A(\u_ps2_keyboard/buffer [4] ), .Z(\u_ps2_keyboard/_0196_ ) );
BUF_X1 \u_ps2_keyboard/_0874_ ( .A(\u_ps2_keyboard/_0100_ ), .Z(\u_ps2_keyboard/_0004_ ) );
BUF_X1 \u_ps2_keyboard/_0875_ ( .A(\u_ps2_keyboard/w_ptr [2] ), .Z(\u_ps2_keyboard/_0448_ ) );
BUF_X1 \u_ps2_keyboard/_0876_ ( .A(\u_ps2_keyboard/w_ptr [1] ), .Z(\u_ps2_keyboard/_0447_ ) );
BUF_X1 \u_ps2_keyboard/_0877_ ( .A(\u_ps2_keyboard/w_ptr [0] ), .Z(\u_ps2_keyboard/_0446_ ) );
BUF_X1 \u_ps2_keyboard/_0878_ ( .A(\u_ps2_keyboard/buffer [0] ), .Z(\u_ps2_keyboard/_0192_ ) );
BUF_X1 \u_ps2_keyboard/_0879_ ( .A(\u_ps2_keyboard/buffer [2] ), .Z(\u_ps2_keyboard/_0194_ ) );
BUF_X1 \u_ps2_keyboard/_0880_ ( .A(\u_ps2_keyboard/buffer [1] ), .Z(\u_ps2_keyboard/_0193_ ) );
BUF_X1 \u_ps2_keyboard/_0881_ ( .A(\u_ps2_keyboard/buffer [3] ), .Z(\u_ps2_keyboard/_0195_ ) );
BUF_X1 \u_ps2_keyboard/_0882_ ( .A(\u_ps2_keyboard/_0174_ ), .Z(\u_ps2_keyboard/_0078_ ) );
BUF_X1 \u_ps2_keyboard/_0883_ ( .A(\u_ps2_keyboard/_0175_ ), .Z(\u_ps2_keyboard/_0079_ ) );
BUF_X1 \u_ps2_keyboard/_0884_ ( .A(\u_ps2_keyboard/_0176_ ), .Z(\u_ps2_keyboard/_0080_ ) );
BUF_X1 \u_ps2_keyboard/_0885_ ( .A(\u_ps2_keyboard/_0177_ ), .Z(\u_ps2_keyboard/_0081_ ) );
BUF_X1 \u_ps2_keyboard/_0886_ ( .A(\u_ps2_keyboard/_0178_ ), .Z(\u_ps2_keyboard/_0082_ ) );
BUF_X1 \u_ps2_keyboard/_0887_ ( .A(\u_ps2_keyboard/_0179_ ), .Z(\u_ps2_keyboard/_0083_ ) );
BUF_X1 \u_ps2_keyboard/_0888_ ( .A(\u_ps2_keyboard/_0180_ ), .Z(\u_ps2_keyboard/_0084_ ) );
BUF_X1 \u_ps2_keyboard/_0889_ ( .A(\u_ps2_keyboard/_0181_ ), .Z(\u_ps2_keyboard/_0085_ ) );
BUF_X1 \u_ps2_keyboard/_0890_ ( .A(\u_ps2_keyboard/_0099_ ), .Z(\u_ps2_keyboard/_0003_ ) );
BUF_X1 \u_ps2_keyboard/_0891_ ( .A(\u_ps2_keyboard/_0166_ ), .Z(\u_ps2_keyboard/_0070_ ) );
BUF_X1 \u_ps2_keyboard/_0892_ ( .A(\u_ps2_keyboard/_0167_ ), .Z(\u_ps2_keyboard/_0071_ ) );
BUF_X1 \u_ps2_keyboard/_0893_ ( .A(\u_ps2_keyboard/_0168_ ), .Z(\u_ps2_keyboard/_0072_ ) );
BUF_X1 \u_ps2_keyboard/_0894_ ( .A(\u_ps2_keyboard/_0169_ ), .Z(\u_ps2_keyboard/_0073_ ) );
BUF_X1 \u_ps2_keyboard/_0895_ ( .A(\u_ps2_keyboard/_0170_ ), .Z(\u_ps2_keyboard/_0074_ ) );
BUF_X1 \u_ps2_keyboard/_0896_ ( .A(\u_ps2_keyboard/_0171_ ), .Z(\u_ps2_keyboard/_0075_ ) );
BUF_X1 \u_ps2_keyboard/_0897_ ( .A(\u_ps2_keyboard/_0172_ ), .Z(\u_ps2_keyboard/_0076_ ) );
BUF_X1 \u_ps2_keyboard/_0898_ ( .A(\u_ps2_keyboard/_0173_ ), .Z(\u_ps2_keyboard/_0077_ ) );
BUF_X1 \u_ps2_keyboard/_0899_ ( .A(\u_ps2_keyboard/_0098_ ), .Z(\u_ps2_keyboard/_0002_ ) );
BUF_X1 \u_ps2_keyboard/_0900_ ( .A(\u_ps2_keyboard/_0097_ ), .Z(\u_ps2_keyboard/_0001_ ) );
BUF_X1 \u_ps2_keyboard/_0901_ ( .A(\u_ps2_keyboard/_0088_ ), .Z(\u_ps2_keyboard/_0184_ ) );
BUF_X1 \u_ps2_keyboard/_0902_ ( .A(\u_ps2_keyboard/_0158_ ), .Z(\u_ps2_keyboard/_0062_ ) );
BUF_X1 \u_ps2_keyboard/_0903_ ( .A(\u_ps2_keyboard/_0159_ ), .Z(\u_ps2_keyboard/_0063_ ) );
BUF_X1 \u_ps2_keyboard/_0904_ ( .A(\u_ps2_keyboard/_0160_ ), .Z(\u_ps2_keyboard/_0064_ ) );
BUF_X1 \u_ps2_keyboard/_0905_ ( .A(\u_ps2_keyboard/_0161_ ), .Z(\u_ps2_keyboard/_0065_ ) );
BUF_X1 \u_ps2_keyboard/_0906_ ( .A(\u_ps2_keyboard/_0162_ ), .Z(\u_ps2_keyboard/_0066_ ) );
BUF_X1 \u_ps2_keyboard/_0907_ ( .A(\u_ps2_keyboard/_0163_ ), .Z(\u_ps2_keyboard/_0067_ ) );
BUF_X1 \u_ps2_keyboard/_0908_ ( .A(\u_ps2_keyboard/_0164_ ), .Z(\u_ps2_keyboard/_0068_ ) );
BUF_X1 \u_ps2_keyboard/_0909_ ( .A(\u_ps2_keyboard/_0165_ ), .Z(\u_ps2_keyboard/_0069_ ) );
BUF_X1 \u_ps2_keyboard/_0910_ ( .A(\u_ps2_keyboard/_0096_ ), .Z(\u_ps2_keyboard/_0000_ ) );
BUF_X1 \u_ps2_keyboard/_0911_ ( .A(\u_ps2_keyboard/_0150_ ), .Z(\u_ps2_keyboard/_0054_ ) );
BUF_X1 \u_ps2_keyboard/_0912_ ( .A(\u_ps2_keyboard/_0151_ ), .Z(\u_ps2_keyboard/_0055_ ) );
BUF_X1 \u_ps2_keyboard/_0913_ ( .A(\u_ps2_keyboard/_0152_ ), .Z(\u_ps2_keyboard/_0056_ ) );
BUF_X1 \u_ps2_keyboard/_0914_ ( .A(\u_ps2_keyboard/_0153_ ), .Z(\u_ps2_keyboard/_0057_ ) );
BUF_X1 \u_ps2_keyboard/_0915_ ( .A(\u_ps2_keyboard/_0154_ ), .Z(\u_ps2_keyboard/_0058_ ) );
BUF_X1 \u_ps2_keyboard/_0916_ ( .A(\u_ps2_keyboard/_0155_ ), .Z(\u_ps2_keyboard/_0059_ ) );
BUF_X1 \u_ps2_keyboard/_0917_ ( .A(\u_ps2_keyboard/_0156_ ), .Z(\u_ps2_keyboard/_0060_ ) );
BUF_X1 \u_ps2_keyboard/_0918_ ( .A(\u_ps2_keyboard/_0157_ ), .Z(\u_ps2_keyboard/_0061_ ) );
BUF_X1 \u_ps2_keyboard/_0919_ ( .A(\u_ps2_keyboard/_0142_ ), .Z(\u_ps2_keyboard/_0046_ ) );
BUF_X1 \u_ps2_keyboard/_0920_ ( .A(\u_ps2_keyboard/_0143_ ), .Z(\u_ps2_keyboard/_0047_ ) );
BUF_X1 \u_ps2_keyboard/_0921_ ( .A(\u_ps2_keyboard/_0144_ ), .Z(\u_ps2_keyboard/_0048_ ) );
BUF_X1 \u_ps2_keyboard/_0922_ ( .A(\u_ps2_keyboard/_0145_ ), .Z(\u_ps2_keyboard/_0049_ ) );
BUF_X1 \u_ps2_keyboard/_0923_ ( .A(\u_ps2_keyboard/_0146_ ), .Z(\u_ps2_keyboard/_0050_ ) );
BUF_X1 \u_ps2_keyboard/_0924_ ( .A(\u_ps2_keyboard/_0147_ ), .Z(\u_ps2_keyboard/_0051_ ) );
BUF_X1 \u_ps2_keyboard/_0925_ ( .A(\u_ps2_keyboard/_0148_ ), .Z(\u_ps2_keyboard/_0052_ ) );
BUF_X1 \u_ps2_keyboard/_0926_ ( .A(\u_ps2_keyboard/_0149_ ), .Z(\u_ps2_keyboard/_0053_ ) );
BUF_X1 \u_ps2_keyboard/_0927_ ( .A(\u_ps2_keyboard/_0115_ ), .Z(\u_ps2_keyboard/_0019_ ) );
BUF_X1 \u_ps2_keyboard/_0928_ ( .A(\u_ps2_keyboard/_0089_ ), .Z(\u_ps2_keyboard/_0185_ ) );
BUF_X1 \u_ps2_keyboard/_0929_ ( .A(\u_ps2_keyboard/_0116_ ), .Z(\u_ps2_keyboard/_0020_ ) );
BUF_X1 \u_ps2_keyboard/_0930_ ( .A(\u_ps2_keyboard/_0090_ ), .Z(\u_ps2_keyboard/_0186_ ) );
BUF_X1 \u_ps2_keyboard/_0931_ ( .A(\u_ps2_keyboard/_0117_ ), .Z(\u_ps2_keyboard/_0021_ ) );
BUF_X1 \u_ps2_keyboard/_0932_ ( .A(_142_ ), .Z(\u_ps2_keyboard/_0428_ ) );
BUF_X1 \u_ps2_keyboard/_0933_ ( .A(\u_ps2_keyboard/_0091_ ), .Z(\u_ps2_keyboard/_0187_ ) );
BUF_X1 \u_ps2_keyboard/_0934_ ( .A(ready ), .Z(\u_ps2_keyboard/_0436_ ) );
BUF_X1 \u_ps2_keyboard/_0935_ ( .A(\u_ps2_keyboard/_0111_ ), .Z(\u_ps2_keyboard/_0015_ ) );
BUF_X1 \u_ps2_keyboard/_0936_ ( .A(\u_ps2_keyboard/_0087_ ), .Z(\u_ps2_keyboard/_0183_ ) );
BUF_X1 \u_ps2_keyboard/_0937_ ( .A(\u_ps2_keyboard/_0112_ ), .Z(\u_ps2_keyboard/_0016_ ) );
BUF_X1 \u_ps2_keyboard/_0938_ ( .A(\u_ps2_keyboard/_0086_ ), .Z(\u_ps2_keyboard/_0182_ ) );
BUF_X1 \u_ps2_keyboard/_0939_ ( .A(\u_ps2_keyboard/_0113_ ), .Z(\u_ps2_keyboard/_0017_ ) );
BUF_X1 \u_ps2_keyboard/_0940_ ( .A(\u_ps2_keyboard/_0134_ ), .Z(\u_ps2_keyboard/_0038_ ) );
BUF_X1 \u_ps2_keyboard/_0941_ ( .A(\u_ps2_keyboard/_0135_ ), .Z(\u_ps2_keyboard/_0039_ ) );
BUF_X1 \u_ps2_keyboard/_0942_ ( .A(\u_ps2_keyboard/_0136_ ), .Z(\u_ps2_keyboard/_0040_ ) );
BUF_X1 \u_ps2_keyboard/_0943_ ( .A(\u_ps2_keyboard/_0137_ ), .Z(\u_ps2_keyboard/_0041_ ) );
BUF_X1 \u_ps2_keyboard/_0944_ ( .A(\u_ps2_keyboard/_0138_ ), .Z(\u_ps2_keyboard/_0042_ ) );
BUF_X1 \u_ps2_keyboard/_0945_ ( .A(\u_ps2_keyboard/_0139_ ), .Z(\u_ps2_keyboard/_0043_ ) );
BUF_X1 \u_ps2_keyboard/_0946_ ( .A(\u_ps2_keyboard/_0140_ ), .Z(\u_ps2_keyboard/_0044_ ) );
BUF_X1 \u_ps2_keyboard/_0947_ ( .A(\u_ps2_keyboard/_0141_ ), .Z(\u_ps2_keyboard/_0045_ ) );
BUF_X1 \u_ps2_keyboard/_0948_ ( .A(\u_ps2_keyboard/_0106_ ), .Z(\u_ps2_keyboard/_0010_ ) );
BUF_X1 \u_ps2_keyboard/_0949_ ( .A(\u_ps2_keyboard/_0092_ ), .Z(\u_ps2_keyboard/_0188_ ) );
BUF_X1 \u_ps2_keyboard/_0950_ ( .A(\u_ps2_keyboard/_0107_ ), .Z(\u_ps2_keyboard/_0011_ ) );
BUF_X1 \u_ps2_keyboard/_0951_ ( .A(\u_ps2_keyboard/_0093_ ), .Z(\u_ps2_keyboard/_0189_ ) );
BUF_X1 \u_ps2_keyboard/_0952_ ( .A(\u_ps2_keyboard/_0108_ ), .Z(\u_ps2_keyboard/_0012_ ) );
BUF_X1 \u_ps2_keyboard/_0953_ ( .A(\u_ps2_keyboard/_0094_ ), .Z(\u_ps2_keyboard/_0190_ ) );
BUF_X1 \u_ps2_keyboard/_0954_ ( .A(\u_ps2_keyboard/_0109_ ), .Z(\u_ps2_keyboard/_0013_ ) );
BUF_X1 \u_ps2_keyboard/_0955_ ( .A(\u_ps2_keyboard/_0126_ ), .Z(\u_ps2_keyboard/_0030_ ) );
BUF_X1 \u_ps2_keyboard/_0956_ ( .A(\u_ps2_keyboard/_0127_ ), .Z(\u_ps2_keyboard/_0031_ ) );
BUF_X1 \u_ps2_keyboard/_0957_ ( .A(\u_ps2_keyboard/_0128_ ), .Z(\u_ps2_keyboard/_0032_ ) );
BUF_X1 \u_ps2_keyboard/_0958_ ( .A(\u_ps2_keyboard/_0129_ ), .Z(\u_ps2_keyboard/_0033_ ) );
BUF_X1 \u_ps2_keyboard/_0959_ ( .A(\u_ps2_keyboard/_0130_ ), .Z(\u_ps2_keyboard/_0034_ ) );
BUF_X1 \u_ps2_keyboard/_0960_ ( .A(\u_ps2_keyboard/_0131_ ), .Z(\u_ps2_keyboard/_0035_ ) );
BUF_X1 \u_ps2_keyboard/_0961_ ( .A(\u_ps2_keyboard/_0132_ ), .Z(\u_ps2_keyboard/_0036_ ) );
BUF_X1 \u_ps2_keyboard/_0962_ ( .A(\u_ps2_keyboard/_0133_ ), .Z(\u_ps2_keyboard/_0037_ ) );
BUF_X1 \u_ps2_keyboard/_0963_ ( .A(\u_ps2_keyboard/_0118_ ), .Z(\u_ps2_keyboard/_0022_ ) );
BUF_X1 \u_ps2_keyboard/_0964_ ( .A(\u_ps2_keyboard/_0119_ ), .Z(\u_ps2_keyboard/_0023_ ) );
BUF_X1 \u_ps2_keyboard/_0965_ ( .A(\u_ps2_keyboard/_0120_ ), .Z(\u_ps2_keyboard/_0024_ ) );
BUF_X1 \u_ps2_keyboard/_0966_ ( .A(\u_ps2_keyboard/_0121_ ), .Z(\u_ps2_keyboard/_0025_ ) );
BUF_X1 \u_ps2_keyboard/_0967_ ( .A(\u_ps2_keyboard/_0122_ ), .Z(\u_ps2_keyboard/_0026_ ) );
BUF_X1 \u_ps2_keyboard/_0968_ ( .A(\u_ps2_keyboard/_0123_ ), .Z(\u_ps2_keyboard/_0027_ ) );
BUF_X1 \u_ps2_keyboard/_0969_ ( .A(\u_ps2_keyboard/_0124_ ), .Z(\u_ps2_keyboard/_0028_ ) );
BUF_X1 \u_ps2_keyboard/_0970_ ( .A(\u_ps2_keyboard/_0125_ ), .Z(\u_ps2_keyboard/_0029_ ) );
BUF_X1 \u_ps2_keyboard/_0971_ ( .A(\u_ps2_keyboard/_0114_ ), .Z(\u_ps2_keyboard/_0018_ ) );
BUF_X1 \u_ps2_keyboard/_0972_ ( .A(overflow ), .Z(\u_ps2_keyboard/_0429_ ) );
BUF_X1 \u_ps2_keyboard/_0973_ ( .A(\u_ps2_keyboard/_0095_ ), .Z(\u_ps2_keyboard/_0191_ ) );
BUF_X1 \u_ps2_keyboard/_0974_ ( .A(\u_ps2_keyboard/_0110_ ), .Z(\u_ps2_keyboard/_0014_ ) );
DFF_X1 \u_ps2_keyboard/_0975_ ( .D(\u_ps2_keyboard/_0070_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[6][0] ), .QN(\u_ps2_keyboard/_0449_ ) );
DFF_X1 \u_ps2_keyboard/_0976_ ( .D(\u_ps2_keyboard/_0071_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[6][1] ), .QN(\u_ps2_keyboard/_0450_ ) );
DFF_X1 \u_ps2_keyboard/_0977_ ( .D(\u_ps2_keyboard/_0072_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[6][2] ), .QN(\u_ps2_keyboard/_0451_ ) );
DFF_X1 \u_ps2_keyboard/_0978_ ( .D(\u_ps2_keyboard/_0073_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[6][3] ), .QN(\u_ps2_keyboard/_0452_ ) );
DFF_X1 \u_ps2_keyboard/_0979_ ( .D(\u_ps2_keyboard/_0074_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[6][4] ), .QN(\u_ps2_keyboard/_0453_ ) );
DFF_X1 \u_ps2_keyboard/_0980_ ( .D(\u_ps2_keyboard/_0075_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[6][5] ), .QN(\u_ps2_keyboard/_0454_ ) );
DFF_X1 \u_ps2_keyboard/_0981_ ( .D(\u_ps2_keyboard/_0076_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[6][6] ), .QN(\u_ps2_keyboard/_0455_ ) );
DFF_X1 \u_ps2_keyboard/_0982_ ( .D(\u_ps2_keyboard/_0077_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[6][7] ), .QN(\u_ps2_keyboard/_0456_ ) );
DFF_X1 \u_ps2_keyboard/_0983_ ( .D(\u_ps2_keyboard/_0015_ ), .CK(clk ), .Q(\u_ps2_keyboard/r_ptr [0] ), .QN(\u_ps2_keyboard/_0091_ ) );
DFF_X1 \u_ps2_keyboard/_0984_ ( .D(\u_ps2_keyboard/_0016_ ), .CK(clk ), .Q(\u_ps2_keyboard/r_ptr [1] ), .QN(\u_ps2_keyboard/_0087_ ) );
DFF_X1 \u_ps2_keyboard/_0985_ ( .D(\u_ps2_keyboard/_0017_ ), .CK(clk ), .Q(\u_ps2_keyboard/r_ptr [2] ), .QN(\u_ps2_keyboard/_0086_ ) );
DFF_X1 \u_ps2_keyboard/_0986_ ( .D(\u_ps2_keyboard/_0022_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[0][0] ), .QN(\u_ps2_keyboard/_0457_ ) );
DFF_X1 \u_ps2_keyboard/_0987_ ( .D(\u_ps2_keyboard/_0023_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[0][1] ), .QN(\u_ps2_keyboard/_0458_ ) );
DFF_X1 \u_ps2_keyboard/_0988_ ( .D(\u_ps2_keyboard/_0024_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[0][2] ), .QN(\u_ps2_keyboard/_0459_ ) );
DFF_X1 \u_ps2_keyboard/_0989_ ( .D(\u_ps2_keyboard/_0025_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[0][3] ), .QN(\u_ps2_keyboard/_0460_ ) );
DFF_X1 \u_ps2_keyboard/_0990_ ( .D(\u_ps2_keyboard/_0026_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[0][4] ), .QN(\u_ps2_keyboard/_0461_ ) );
DFF_X1 \u_ps2_keyboard/_0991_ ( .D(\u_ps2_keyboard/_0027_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[0][5] ), .QN(\u_ps2_keyboard/_0462_ ) );
DFF_X1 \u_ps2_keyboard/_0992_ ( .D(\u_ps2_keyboard/_0028_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[0][6] ), .QN(\u_ps2_keyboard/_0463_ ) );
DFF_X1 \u_ps2_keyboard/_0993_ ( .D(\u_ps2_keyboard/_0029_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[0][7] ), .QN(\u_ps2_keyboard/_0464_ ) );
DFF_X1 \u_ps2_keyboard/_0994_ ( .D(\u_ps2_keyboard/_0030_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[1][0] ), .QN(\u_ps2_keyboard/_0465_ ) );
DFF_X1 \u_ps2_keyboard/_0995_ ( .D(\u_ps2_keyboard/_0031_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[1][1] ), .QN(\u_ps2_keyboard/_0466_ ) );
DFF_X1 \u_ps2_keyboard/_0996_ ( .D(\u_ps2_keyboard/_0032_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[1][2] ), .QN(\u_ps2_keyboard/_0467_ ) );
DFF_X1 \u_ps2_keyboard/_0997_ ( .D(\u_ps2_keyboard/_0033_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[1][3] ), .QN(\u_ps2_keyboard/_0468_ ) );
DFF_X1 \u_ps2_keyboard/_0998_ ( .D(\u_ps2_keyboard/_0034_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[1][4] ), .QN(\u_ps2_keyboard/_0469_ ) );
DFF_X1 \u_ps2_keyboard/_0999_ ( .D(\u_ps2_keyboard/_0035_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[1][5] ), .QN(\u_ps2_keyboard/_0470_ ) );
DFF_X1 \u_ps2_keyboard/_1000_ ( .D(\u_ps2_keyboard/_0036_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[1][6] ), .QN(\u_ps2_keyboard/_0471_ ) );
DFF_X1 \u_ps2_keyboard/_1001_ ( .D(\u_ps2_keyboard/_0037_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[1][7] ), .QN(\u_ps2_keyboard/_0472_ ) );
DFF_X1 \u_ps2_keyboard/_1002_ ( .D(\u_ps2_keyboard/_0046_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[3][0] ), .QN(\u_ps2_keyboard/_0473_ ) );
DFF_X1 \u_ps2_keyboard/_1003_ ( .D(\u_ps2_keyboard/_0047_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[3][1] ), .QN(\u_ps2_keyboard/_0474_ ) );
DFF_X1 \u_ps2_keyboard/_1004_ ( .D(\u_ps2_keyboard/_0048_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[3][2] ), .QN(\u_ps2_keyboard/_0475_ ) );
DFF_X1 \u_ps2_keyboard/_1005_ ( .D(\u_ps2_keyboard/_0049_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[3][3] ), .QN(\u_ps2_keyboard/_0476_ ) );
DFF_X1 \u_ps2_keyboard/_1006_ ( .D(\u_ps2_keyboard/_0050_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[3][4] ), .QN(\u_ps2_keyboard/_0477_ ) );
DFF_X1 \u_ps2_keyboard/_1007_ ( .D(\u_ps2_keyboard/_0051_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[3][5] ), .QN(\u_ps2_keyboard/_0478_ ) );
DFF_X1 \u_ps2_keyboard/_1008_ ( .D(\u_ps2_keyboard/_0052_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[3][6] ), .QN(\u_ps2_keyboard/_0479_ ) );
DFF_X1 \u_ps2_keyboard/_1009_ ( .D(\u_ps2_keyboard/_0053_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[3][7] ), .QN(\u_ps2_keyboard/_0480_ ) );
DFF_X1 \u_ps2_keyboard/_1010_ ( .D(\u_ps2_keyboard/_0054_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[4][0] ), .QN(\u_ps2_keyboard/_0481_ ) );
DFF_X1 \u_ps2_keyboard/_1011_ ( .D(\u_ps2_keyboard/_0055_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[4][1] ), .QN(\u_ps2_keyboard/_0482_ ) );
DFF_X1 \u_ps2_keyboard/_1012_ ( .D(\u_ps2_keyboard/_0056_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[4][2] ), .QN(\u_ps2_keyboard/_0483_ ) );
DFF_X1 \u_ps2_keyboard/_1013_ ( .D(\u_ps2_keyboard/_0057_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[4][3] ), .QN(\u_ps2_keyboard/_0484_ ) );
DFF_X1 \u_ps2_keyboard/_1014_ ( .D(\u_ps2_keyboard/_0058_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[4][4] ), .QN(\u_ps2_keyboard/_0485_ ) );
DFF_X1 \u_ps2_keyboard/_1015_ ( .D(\u_ps2_keyboard/_0059_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[4][5] ), .QN(\u_ps2_keyboard/_0486_ ) );
DFF_X1 \u_ps2_keyboard/_1016_ ( .D(\u_ps2_keyboard/_0060_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[4][6] ), .QN(\u_ps2_keyboard/_0487_ ) );
DFF_X1 \u_ps2_keyboard/_1017_ ( .D(\u_ps2_keyboard/_0061_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[4][7] ), .QN(\u_ps2_keyboard/_0488_ ) );
DFF_X1 \u_ps2_keyboard/_1018_ ( .D(\u_ps2_keyboard/_0038_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[2][0] ), .QN(\u_ps2_keyboard/_0489_ ) );
DFF_X1 \u_ps2_keyboard/_1019_ ( .D(\u_ps2_keyboard/_0039_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[2][1] ), .QN(\u_ps2_keyboard/_0490_ ) );
DFF_X1 \u_ps2_keyboard/_1020_ ( .D(\u_ps2_keyboard/_0040_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[2][2] ), .QN(\u_ps2_keyboard/_0491_ ) );
DFF_X1 \u_ps2_keyboard/_1021_ ( .D(\u_ps2_keyboard/_0041_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[2][3] ), .QN(\u_ps2_keyboard/_0492_ ) );
DFF_X1 \u_ps2_keyboard/_1022_ ( .D(\u_ps2_keyboard/_0042_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[2][4] ), .QN(\u_ps2_keyboard/_0493_ ) );
DFF_X1 \u_ps2_keyboard/_1023_ ( .D(\u_ps2_keyboard/_0043_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[2][5] ), .QN(\u_ps2_keyboard/_0494_ ) );
DFF_X1 \u_ps2_keyboard/_1024_ ( .D(\u_ps2_keyboard/_0044_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[2][6] ), .QN(\u_ps2_keyboard/_0495_ ) );
DFF_X1 \u_ps2_keyboard/_1025_ ( .D(\u_ps2_keyboard/_0045_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[2][7] ), .QN(\u_ps2_keyboard/_0496_ ) );
DFF_X1 \u_ps2_keyboard/_1026_ ( .D(\u_ps2_keyboard/_0078_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[7][0] ), .QN(\u_ps2_keyboard/_0497_ ) );
DFF_X1 \u_ps2_keyboard/_1027_ ( .D(\u_ps2_keyboard/_0079_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[7][1] ), .QN(\u_ps2_keyboard/_0498_ ) );
DFF_X1 \u_ps2_keyboard/_1028_ ( .D(\u_ps2_keyboard/_0080_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[7][2] ), .QN(\u_ps2_keyboard/_0499_ ) );
DFF_X1 \u_ps2_keyboard/_1029_ ( .D(\u_ps2_keyboard/_0081_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[7][3] ), .QN(\u_ps2_keyboard/_0500_ ) );
DFF_X1 \u_ps2_keyboard/_1030_ ( .D(\u_ps2_keyboard/_0082_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[7][4] ), .QN(\u_ps2_keyboard/_0501_ ) );
DFF_X1 \u_ps2_keyboard/_1031_ ( .D(\u_ps2_keyboard/_0083_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[7][5] ), .QN(\u_ps2_keyboard/_0502_ ) );
DFF_X1 \u_ps2_keyboard/_1032_ ( .D(\u_ps2_keyboard/_0084_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[7][6] ), .QN(\u_ps2_keyboard/_0503_ ) );
DFF_X1 \u_ps2_keyboard/_1033_ ( .D(\u_ps2_keyboard/_0085_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[7][7] ), .QN(\u_ps2_keyboard/_0504_ ) );
DFF_X1 \u_ps2_keyboard/_1034_ ( .D(\u_ps2_keyboard/_0018_ ), .CK(clk ), .Q(ready ), .QN(\u_ps2_keyboard/_0505_ ) );
DFF_X1 \u_ps2_keyboard/_1035_ ( .D(\u_ps2_keyboard/_0062_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[5][0] ), .QN(\u_ps2_keyboard/_0506_ ) );
DFF_X1 \u_ps2_keyboard/_1036_ ( .D(\u_ps2_keyboard/_0063_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[5][1] ), .QN(\u_ps2_keyboard/_0507_ ) );
DFF_X1 \u_ps2_keyboard/_1037_ ( .D(\u_ps2_keyboard/_0064_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[5][2] ), .QN(\u_ps2_keyboard/_0508_ ) );
DFF_X1 \u_ps2_keyboard/_1038_ ( .D(\u_ps2_keyboard/_0065_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[5][3] ), .QN(\u_ps2_keyboard/_0509_ ) );
DFF_X1 \u_ps2_keyboard/_1039_ ( .D(\u_ps2_keyboard/_0066_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[5][4] ), .QN(\u_ps2_keyboard/_0510_ ) );
DFF_X1 \u_ps2_keyboard/_1040_ ( .D(\u_ps2_keyboard/_0067_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[5][5] ), .QN(\u_ps2_keyboard/_0511_ ) );
DFF_X1 \u_ps2_keyboard/_1041_ ( .D(\u_ps2_keyboard/_0068_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[5][6] ), .QN(\u_ps2_keyboard/_0512_ ) );
DFF_X1 \u_ps2_keyboard/_1042_ ( .D(\u_ps2_keyboard/_0069_ ), .CK(clk ), .Q(\u_ps2_keyboard/fifo[5][7] ), .QN(\u_ps2_keyboard/_0513_ ) );
DFF_X1 \u_ps2_keyboard/_1043_ ( .D(\u_ps2_keyboard/_0014_ ), .CK(clk ), .Q(overflow ), .QN(\u_ps2_keyboard/_0095_ ) );
DFF_X1 \u_ps2_keyboard/_1044_ ( .D(\u_ps2_keyboard/_0010_ ), .CK(clk ), .Q(\u_ps2_keyboard/count [0] ), .QN(\u_ps2_keyboard/_0514_ ) );
DFF_X1 \u_ps2_keyboard/_1045_ ( .D(\u_ps2_keyboard/_0011_ ), .CK(clk ), .Q(\u_ps2_keyboard/count [1] ), .QN(\u_ps2_keyboard/_0092_ ) );
DFF_X1 \u_ps2_keyboard/_1046_ ( .D(\u_ps2_keyboard/_0012_ ), .CK(clk ), .Q(\u_ps2_keyboard/count [2] ), .QN(\u_ps2_keyboard/_0093_ ) );
DFF_X1 \u_ps2_keyboard/_1047_ ( .D(\u_ps2_keyboard/_0013_ ), .CK(clk ), .Q(\u_ps2_keyboard/count [3] ), .QN(\u_ps2_keyboard/_0094_ ) );
DFF_X1 \u_ps2_keyboard/_1048_ ( .D(\u_ps2_keyboard/_0019_ ), .CK(clk ), .Q(\u_ps2_keyboard/w_ptr [0] ), .QN(\u_ps2_keyboard/_0088_ ) );
DFF_X1 \u_ps2_keyboard/_1049_ ( .D(\u_ps2_keyboard/_0020_ ), .CK(clk ), .Q(\u_ps2_keyboard/w_ptr [1] ), .QN(\u_ps2_keyboard/_0089_ ) );
DFF_X1 \u_ps2_keyboard/_1050_ ( .D(\u_ps2_keyboard/_0021_ ), .CK(clk ), .Q(\u_ps2_keyboard/w_ptr [2] ), .QN(\u_ps2_keyboard/_0090_ ) );
DFF_X1 \u_ps2_keyboard/_1051_ ( .D(\u_ps2_keyboard/_0000_ ), .CK(clk ), .Q(\u_ps2_keyboard/buffer [0] ), .QN(\u_ps2_keyboard/_0515_ ) );
DFF_X1 \u_ps2_keyboard/_1052_ ( .D(\u_ps2_keyboard/_0001_ ), .CK(clk ), .Q(\u_ps2_keyboard/buffer [1] ), .QN(\u_ps2_keyboard/_0516_ ) );
DFF_X1 \u_ps2_keyboard/_1053_ ( .D(\u_ps2_keyboard/_0002_ ), .CK(clk ), .Q(\u_ps2_keyboard/buffer [2] ), .QN(\u_ps2_keyboard/_0517_ ) );
DFF_X1 \u_ps2_keyboard/_1054_ ( .D(\u_ps2_keyboard/_0003_ ), .CK(clk ), .Q(\u_ps2_keyboard/buffer [3] ), .QN(\u_ps2_keyboard/_0518_ ) );
DFF_X1 \u_ps2_keyboard/_1055_ ( .D(\u_ps2_keyboard/_0004_ ), .CK(clk ), .Q(\u_ps2_keyboard/buffer [4] ), .QN(\u_ps2_keyboard/_0519_ ) );
DFF_X1 \u_ps2_keyboard/_1056_ ( .D(\u_ps2_keyboard/_0005_ ), .CK(clk ), .Q(\u_ps2_keyboard/buffer [5] ), .QN(\u_ps2_keyboard/_0520_ ) );
DFF_X1 \u_ps2_keyboard/_1057_ ( .D(\u_ps2_keyboard/_0006_ ), .CK(clk ), .Q(\u_ps2_keyboard/buffer [6] ), .QN(\u_ps2_keyboard/_0521_ ) );
DFF_X1 \u_ps2_keyboard/_1058_ ( .D(\u_ps2_keyboard/_0007_ ), .CK(clk ), .Q(\u_ps2_keyboard/buffer [7] ), .QN(\u_ps2_keyboard/_0522_ ) );
DFF_X1 \u_ps2_keyboard/_1059_ ( .D(\u_ps2_keyboard/_0008_ ), .CK(clk ), .Q(\u_ps2_keyboard/buffer [8] ), .QN(\u_ps2_keyboard/_0523_ ) );
DFF_X1 \u_ps2_keyboard/_1060_ ( .D(\u_ps2_keyboard/_0009_ ), .CK(clk ), .Q(\u_ps2_keyboard/buffer [9] ), .QN(\u_ps2_keyboard/_0524_ ) );
DFF_X1 \u_ps2_keyboard/_1061_ ( .D(ps2_clk ), .CK(clk ), .Q(\u_ps2_keyboard/ps2_clk_sync [0] ), .QN(\u_ps2_keyboard/_0525_ ) );
DFF_X1 \u_ps2_keyboard/_1062_ ( .D(\u_ps2_keyboard/ps2_clk_sync [0] ), .CK(clk ), .Q(\u_ps2_keyboard/ps2_clk_sync [1] ), .QN(\u_ps2_keyboard/_0526_ ) );
DFF_X1 \u_ps2_keyboard/_1063_ ( .D(\u_ps2_keyboard/ps2_clk_sync [1] ), .CK(clk ), .Q(\u_ps2_keyboard/ps2_clk_sync [2] ), .QN(\u_ps2_keyboard/_0527_ ) );
NOR2_X4 \u_rom/_050_ ( .A1(\u_rom/_048_ ), .A2(\u_rom/_047_ ), .ZN(\u_rom/_007_ ) );
INV_X16 \u_rom/_051_ ( .A(\u_rom/_046_ ), .ZN(\u_rom/_008_ ) );
AND3_X4 \u_rom/_052_ ( .A1(\u_rom/_007_ ), .A2(\u_rom/_008_ ), .A3(\u_rom/_045_ ), .ZN(\u_rom/_009_ ) );
INV_X32 \u_rom/_053_ ( .A(\u_rom/_043_ ), .ZN(\u_rom/_010_ ) );
NOR2_X4 \u_rom/_054_ ( .A1(\u_rom/_010_ ), .A2(\u_rom/_044_ ), .ZN(\u_rom/_011_ ) );
INV_X32 \u_rom/_055_ ( .A(\u_rom/_042_ ), .ZN(\u_rom/_012_ ) );
AND3_X4 \u_rom/_056_ ( .A1(\u_rom/_011_ ), .A2(\u_rom/_012_ ), .A3(\u_rom/_041_ ), .ZN(\u_rom/_013_ ) );
NOR2_X4 \u_rom/_057_ ( .A1(\u_rom/_012_ ), .A2(\u_rom/_041_ ), .ZN(\u_rom/_014_ ) );
AND2_X1 \u_rom/_058_ ( .A1(\u_rom/_011_ ), .A2(\u_rom/_014_ ), .ZN(\u_rom/_015_ ) );
OAI21_X1 \u_rom/_059_ ( .A(\u_rom/_009_ ), .B1(\u_rom/_013_ ), .B2(\u_rom/_015_ ), .ZN(\u_rom/_016_ ) );
NOR2_X2 \u_rom/_060_ ( .A1(\u_rom/_008_ ), .A2(\u_rom/_047_ ), .ZN(\u_rom/_017_ ) );
NOR2_X4 \u_rom/_061_ ( .A1(\u_rom/_045_ ), .A2(\u_rom/_048_ ), .ZN(\u_rom/_018_ ) );
AND2_X1 \u_rom/_062_ ( .A1(\u_rom/_017_ ), .A2(\u_rom/_018_ ), .ZN(\u_rom/_019_ ) );
AND3_X1 \u_rom/_063_ ( .A1(\u_rom/_019_ ), .A2(\u_rom/_043_ ), .A3(\u_rom/_014_ ), .ZN(\u_rom/_020_ ) );
AND3_X2 \u_rom/_064_ ( .A1(\u_rom/_018_ ), .A2(\u_rom/_008_ ), .A3(\u_rom/_047_ ), .ZN(\u_rom/_021_ ) );
AND3_X2 \u_rom/_065_ ( .A1(\u_rom/_021_ ), .A2(\u_rom/_011_ ), .A3(\u_rom/_014_ ), .ZN(\u_rom/_022_ ) );
AND2_X4 \u_rom/_066_ ( .A1(\u_rom/_044_ ), .A2(\u_rom/_043_ ), .ZN(\u_rom/_023_ ) );
AND3_X1 \u_rom/_067_ ( .A1(\u_rom/_023_ ), .A2(\u_rom/_012_ ), .A3(\u_rom/_041_ ), .ZN(\u_rom/_024_ ) );
AND2_X4 \u_rom/_068_ ( .A1(\u_rom/_046_ ), .A2(\u_rom/_045_ ), .ZN(\u_rom/_025_ ) );
AND2_X1 \u_rom/_069_ ( .A1(\u_rom/_025_ ), .A2(\u_rom/_007_ ), .ZN(\u_rom/_026_ ) );
AND2_X2 \u_rom/_070_ ( .A1(\u_rom/_024_ ), .A2(\u_rom/_026_ ), .ZN(\u_rom/_027_ ) );
NOR3_X1 \u_rom/_071_ ( .A1(\u_rom/_020_ ), .A2(\u_rom/_022_ ), .A3(\u_rom/_027_ ), .ZN(\u_rom/_028_ ) );
AND3_X2 \u_rom/_072_ ( .A1(\u_rom/_009_ ), .A2(\u_rom/_014_ ), .A3(\u_rom/_023_ ), .ZN(\u_rom/_029_ ) );
AND4_X2 \u_rom/_073_ ( .A1(\u_rom/_007_ ), .A2(\u_rom/_011_ ), .A3(\u_rom/_014_ ), .A4(\u_rom/_025_ ), .ZN(\u_rom/_030_ ) );
AND4_X1 \u_rom/_074_ ( .A1(\u_rom/_018_ ), .A2(\u_rom/_017_ ), .A3(\u_rom/_011_ ), .A4(\u_rom/_014_ ), .ZN(\u_rom/_031_ ) );
OR4_X4 \u_rom/_075_ ( .A1(\u_rom/_027_ ), .A2(\u_rom/_029_ ), .A3(\u_rom/_030_ ), .A4(\u_rom/_031_ ), .ZN(\u_rom/_001_ ) );
AND2_X1 \u_rom/_076_ ( .A1(\u_rom/_014_ ), .A2(\u_rom/_023_ ), .ZN(\u_rom/_032_ ) );
NOR2_X2 \u_rom/_077_ ( .A1(\u_rom/_013_ ), .A2(\u_rom/_032_ ), .ZN(\u_rom/_033_ ) );
INV_X1 \u_rom/_078_ ( .A(\u_rom/_019_ ), .ZN(\u_rom/_034_ ) );
NOR2_X2 \u_rom/_079_ ( .A1(\u_rom/_033_ ), .A2(\u_rom/_034_ ), .ZN(\u_rom/_035_ ) );
AND4_X1 \u_rom/_080_ ( .A1(\u_rom/_007_ ), .A2(\u_rom/_014_ ), .A3(\u_rom/_023_ ), .A4(\u_rom/_025_ ), .ZN(\u_rom/_036_ ) );
OR2_X2 \u_rom/_081_ ( .A1(\u_rom/_036_ ), .A2(\u_rom/_022_ ), .ZN(\u_rom/_003_ ) );
NOR3_X4 \u_rom/_082_ ( .A1(\u_rom/_001_ ), .A2(\u_rom/_035_ ), .A3(\u_rom/_003_ ), .ZN(\u_rom/_037_ ) );
INV_X1 \u_rom/_083_ ( .A(\u_rom/_037_ ), .ZN(\u_rom/_038_ ) );
AND2_X1 \u_rom/_084_ ( .A1(\u_rom/_013_ ), .A2(\u_rom/_021_ ), .ZN(\u_rom/_039_ ) );
OAI211_X2 \u_rom/_085_ ( .A(\u_rom/_016_ ), .B(\u_rom/_028_ ), .C1(\u_rom/_038_ ), .C2(\u_rom/_039_ ), .ZN(\u_rom/_000_ ) );
OR3_X1 \u_rom/_086_ ( .A1(\u_rom/_035_ ), .A2(\u_rom/_027_ ), .A3(\u_rom/_030_ ), .ZN(\u_rom/_002_ ) );
AND2_X1 \u_rom/_087_ ( .A1(\u_rom/_013_ ), .A2(\u_rom/_009_ ), .ZN(\u_rom/_004_ ) );
AOI21_X1 \u_rom/_088_ ( .A(\u_rom/_039_ ), .B1(\u_rom/_015_ ), .B2(\u_rom/_009_ ), .ZN(\u_rom/_040_ ) );
AND2_X2 \u_rom/_089_ ( .A1(\u_rom/_037_ ), .A2(\u_rom/_040_ ), .ZN(\u_rom/_006_ ) );
INV_X1 \u_rom/_090_ ( .A(\u_rom/_006_ ), .ZN(\u_rom/_005_ ) );
LOGIC0_X1 \u_rom/_091_ ( .Z(\u_rom/_049_ ) );
BUF_X1 \u_rom/_092_ ( .A(\u_rom/_049_ ), .Z(\ascii_code [7] ) );
BUF_X1 \u_rom/_093_ ( .A(\scan_code_buf [1] ), .Z(\u_rom/_042_ ) );
BUF_X1 \u_rom/_094_ ( .A(\scan_code_buf [0] ), .Z(\u_rom/_041_ ) );
BUF_X1 \u_rom/_095_ ( .A(\scan_code_buf [3] ), .Z(\u_rom/_044_ ) );
BUF_X1 \u_rom/_096_ ( .A(\scan_code_buf [2] ), .Z(\u_rom/_043_ ) );
BUF_X1 \u_rom/_097_ ( .A(\scan_code_buf [5] ), .Z(\u_rom/_046_ ) );
BUF_X1 \u_rom/_098_ ( .A(\scan_code_buf [4] ), .Z(\u_rom/_045_ ) );
BUF_X1 \u_rom/_099_ ( .A(\scan_code_buf [7] ), .Z(\u_rom/_048_ ) );
BUF_X1 \u_rom/_100_ ( .A(\scan_code_buf [6] ), .Z(\u_rom/_047_ ) );
BUF_X1 \u_rom/_101_ ( .A(\u_rom/_000_ ), .Z(\ascii_code [0] ) );
BUF_X1 \u_rom/_102_ ( .A(\u_rom/_001_ ), .Z(\ascii_code [1] ) );
BUF_X1 \u_rom/_103_ ( .A(\u_rom/_002_ ), .Z(\ascii_code [2] ) );
BUF_X1 \u_rom/_104_ ( .A(\u_rom/_003_ ), .Z(\ascii_code [3] ) );
BUF_X1 \u_rom/_105_ ( .A(\u_rom/_004_ ), .Z(\ascii_code [4] ) );
BUF_X1 \u_rom/_106_ ( .A(\u_rom/_005_ ), .Z(\ascii_code [5] ) );
BUF_X1 \u_rom/_107_ ( .A(\u_rom/_006_ ), .Z(\ascii_code [6] ) );
NOR2_X4 \u_scan_code_h/_43_ ( .A1(\u_scan_code_h/_01_ ), .A2(\u_scan_code_h/_00_ ), .ZN(\u_scan_code_h/_05_ ) );
INV_X2 \u_scan_code_h/_44_ ( .A(\u_scan_code_h/_05_ ), .ZN(\u_scan_code_h/_06_ ) );
INV_X4 \u_scan_code_h/_45_ ( .A(\u_scan_code_h/_02_ ), .ZN(\u_scan_code_h/_07_ ) );
NOR2_X2 \u_scan_code_h/_46_ ( .A1(\u_scan_code_h/_07_ ), .A2(\u_scan_code_h/_03_ ), .ZN(\u_scan_code_h/_08_ ) );
INV_X16 \u_scan_code_h/_47_ ( .A(\u_scan_code_h/_03_ ), .ZN(\u_scan_code_h/_09_ ) );
NOR2_X2 \u_scan_code_h/_48_ ( .A1(\u_scan_code_h/_09_ ), .A2(\u_scan_code_h/_02_ ), .ZN(\u_scan_code_h/_10_ ) );
OR3_X4 \u_scan_code_h/_49_ ( .A1(\u_scan_code_h/_06_ ), .A2(\u_scan_code_h/_08_ ), .A3(\u_scan_code_h/_10_ ), .ZN(\u_scan_code_h/_11_ ) );
INV_X32 \u_scan_code_h/_50_ ( .A(\u_scan_code_h/_00_ ), .ZN(\u_scan_code_h/_12_ ) );
NOR2_X2 \u_scan_code_h/_51_ ( .A1(\u_scan_code_h/_12_ ), .A2(\u_scan_code_h/_01_ ), .ZN(\u_scan_code_h/_13_ ) );
NOR2_X4 \u_scan_code_h/_52_ ( .A1(\u_scan_code_h/_03_ ), .A2(\u_scan_code_h/_02_ ), .ZN(\u_scan_code_h/_14_ ) );
AND2_X1 \u_scan_code_h/_53_ ( .A1(\u_scan_code_h/_13_ ), .A2(\u_scan_code_h/_14_ ), .ZN(\u_scan_code_h/_15_ ) );
INV_X1 \u_scan_code_h/_54_ ( .A(\u_scan_code_h/_15_ ), .ZN(\u_scan_code_h/_16_ ) );
INV_X1 \u_scan_code_h/_55_ ( .A(\u_scan_code_h/_04_ ), .ZN(\u_scan_code_h/_17_ ) );
AND2_X4 \u_scan_code_h/_56_ ( .A1(\u_scan_code_h/_01_ ), .A2(\u_scan_code_h/_00_ ), .ZN(\u_scan_code_h/_18_ ) );
AOI21_X1 \u_scan_code_h/_57_ ( .A(\u_scan_code_h/_17_ ), .B1(\u_scan_code_h/_08_ ), .B2(\u_scan_code_h/_18_ ), .ZN(\u_scan_code_h/_19_ ) );
NAND3_X1 \u_scan_code_h/_58_ ( .A1(\u_scan_code_h/_11_ ), .A2(\u_scan_code_h/_16_ ), .A3(\u_scan_code_h/_19_ ), .ZN(\u_scan_code_h/_35_ ) );
NAND2_X1 \u_scan_code_h/_59_ ( .A1(\u_scan_code_h/_06_ ), .A2(\u_scan_code_h/_14_ ), .ZN(\u_scan_code_h/_20_ ) );
AND2_X2 \u_scan_code_h/_60_ ( .A1(\u_scan_code_h/_03_ ), .A2(\u_scan_code_h/_02_ ), .ZN(\u_scan_code_h/_21_ ) );
NAND2_X1 \u_scan_code_h/_61_ ( .A1(\u_scan_code_h/_13_ ), .A2(\u_scan_code_h/_21_ ), .ZN(\u_scan_code_h/_22_ ) );
NAND3_X1 \u_scan_code_h/_62_ ( .A1(\u_scan_code_h/_19_ ), .A2(\u_scan_code_h/_20_ ), .A3(\u_scan_code_h/_22_ ), .ZN(\u_scan_code_h/_36_ ) );
NOR3_X1 \u_scan_code_h/_63_ ( .A1(\u_scan_code_h/_07_ ), .A2(\u_scan_code_h/_03_ ), .A3(\u_scan_code_h/_01_ ), .ZN(\u_scan_code_h/_23_ ) );
AOI21_X1 \u_scan_code_h/_64_ ( .A(\u_scan_code_h/_23_ ), .B1(\u_scan_code_h/_08_ ), .B2(\u_scan_code_h/_18_ ), .ZN(\u_scan_code_h/_24_ ) );
NAND3_X1 \u_scan_code_h/_65_ ( .A1(\u_scan_code_h/_09_ ), .A2(\u_scan_code_h/_07_ ), .A3(\u_scan_code_h/_00_ ), .ZN(\u_scan_code_h/_25_ ) );
NAND2_X1 \u_scan_code_h/_66_ ( .A1(\u_scan_code_h/_13_ ), .A2(\u_scan_code_h/_10_ ), .ZN(\u_scan_code_h/_26_ ) );
NAND4_X1 \u_scan_code_h/_67_ ( .A1(\u_scan_code_h/_24_ ), .A2(\u_scan_code_h/_04_ ), .A3(\u_scan_code_h/_25_ ), .A4(\u_scan_code_h/_26_ ), .ZN(\u_scan_code_h/_37_ ) );
NAND3_X1 \u_scan_code_h/_68_ ( .A1(\u_scan_code_h/_10_ ), .A2(\u_scan_code_h/_01_ ), .A3(\u_scan_code_h/_12_ ), .ZN(\u_scan_code_h/_27_ ) );
AOI22_X1 \u_scan_code_h/_69_ ( .A1(\u_scan_code_h/_08_ ), .A2(\u_scan_code_h/_05_ ), .B1(\u_scan_code_h/_18_ ), .B2(\u_scan_code_h/_21_ ), .ZN(\u_scan_code_h/_28_ ) );
NAND4_X1 \u_scan_code_h/_70_ ( .A1(\u_scan_code_h/_16_ ), .A2(\u_scan_code_h/_19_ ), .A3(\u_scan_code_h/_27_ ), .A4(\u_scan_code_h/_28_ ), .ZN(\u_scan_code_h/_38_ ) );
OAI21_X1 \u_scan_code_h/_71_ ( .A(\u_scan_code_h/_21_ ), .B1(\u_scan_code_h/_01_ ), .B2(\u_scan_code_h/_12_ ), .ZN(\u_scan_code_h/_29_ ) );
NAND3_X1 \u_scan_code_h/_72_ ( .A1(\u_scan_code_h/_14_ ), .A2(\u_scan_code_h/_01_ ), .A3(\u_scan_code_h/_12_ ), .ZN(\u_scan_code_h/_30_ ) );
NAND3_X1 \u_scan_code_h/_73_ ( .A1(\u_scan_code_h/_29_ ), .A2(\u_scan_code_h/_30_ ), .A3(\u_scan_code_h/_04_ ), .ZN(\u_scan_code_h/_39_ ) );
AND2_X1 \u_scan_code_h/_74_ ( .A1(\u_scan_code_h/_12_ ), .A2(\u_scan_code_h/_01_ ), .ZN(\u_scan_code_h/_31_ ) );
OAI21_X1 \u_scan_code_h/_75_ ( .A(\u_scan_code_h/_08_ ), .B1(\u_scan_code_h/_31_ ), .B2(\u_scan_code_h/_13_ ), .ZN(\u_scan_code_h/_32_ ) );
NAND2_X1 \u_scan_code_h/_76_ ( .A1(\u_scan_code_h/_10_ ), .A2(\u_scan_code_h/_18_ ), .ZN(\u_scan_code_h/_33_ ) );
NAND4_X1 \u_scan_code_h/_77_ ( .A1(\u_scan_code_h/_32_ ), .A2(\u_scan_code_h/_04_ ), .A3(\u_scan_code_h/_29_ ), .A4(\u_scan_code_h/_33_ ), .ZN(\u_scan_code_h/_40_ ) );
AOI22_X1 \u_scan_code_h/_78_ ( .A1(\u_scan_code_h/_14_ ), .A2(\u_scan_code_h/_13_ ), .B1(\u_scan_code_h/_08_ ), .B2(\u_scan_code_h/_05_ ), .ZN(\u_scan_code_h/_34_ ) );
NAND4_X1 \u_scan_code_h/_79_ ( .A1(\u_scan_code_h/_34_ ), .A2(\u_scan_code_h/_04_ ), .A3(\u_scan_code_h/_22_ ), .A4(\u_scan_code_h/_33_ ), .ZN(\u_scan_code_h/_41_ ) );
LOGIC1_X1 \u_scan_code_h/_80_ ( .Z(\u_scan_code_h/_42_ ) );
BUF_X1 \u_scan_code_h/_81_ ( .A(\u_scan_code_h/_42_ ), .Z(\scan_code_seg [8] ) );
BUF_X1 \u_scan_code_h/_82_ ( .A(\scan_code_buf [7] ), .Z(\u_scan_code_h/_03_ ) );
BUF_X1 \u_scan_code_h/_83_ ( .A(\scan_code_buf [6] ), .Z(\u_scan_code_h/_02_ ) );
BUF_X1 \u_scan_code_h/_84_ ( .A(\scan_code_buf [5] ), .Z(\u_scan_code_h/_01_ ) );
BUF_X1 \u_scan_code_h/_85_ ( .A(\scan_code_buf [4] ), .Z(\u_scan_code_h/_00_ ) );
BUF_X1 \u_scan_code_h/_86_ ( .A(display_en ), .Z(\u_scan_code_h/_04_ ) );
BUF_X1 \u_scan_code_h/_87_ ( .A(\u_scan_code_h/_35_ ), .Z(\scan_code_seg [9] ) );
BUF_X1 \u_scan_code_h/_88_ ( .A(\u_scan_code_h/_36_ ), .Z(\scan_code_seg [10] ) );
BUF_X1 \u_scan_code_h/_89_ ( .A(\u_scan_code_h/_37_ ), .Z(\scan_code_seg [11] ) );
BUF_X1 \u_scan_code_h/_90_ ( .A(\u_scan_code_h/_38_ ), .Z(\scan_code_seg [12] ) );
BUF_X1 \u_scan_code_h/_91_ ( .A(\u_scan_code_h/_39_ ), .Z(\scan_code_seg [13] ) );
BUF_X1 \u_scan_code_h/_92_ ( .A(\u_scan_code_h/_40_ ), .Z(\scan_code_seg [14] ) );
BUF_X1 \u_scan_code_h/_93_ ( .A(\u_scan_code_h/_41_ ), .Z(\scan_code_seg [15] ) );
NOR2_X4 \u_scan_code_l/_43_ ( .A1(\u_scan_code_l/_01_ ), .A2(\u_scan_code_l/_00_ ), .ZN(\u_scan_code_l/_05_ ) );
INV_X2 \u_scan_code_l/_44_ ( .A(\u_scan_code_l/_05_ ), .ZN(\u_scan_code_l/_06_ ) );
INV_X4 \u_scan_code_l/_45_ ( .A(\u_scan_code_l/_02_ ), .ZN(\u_scan_code_l/_07_ ) );
NOR2_X2 \u_scan_code_l/_46_ ( .A1(\u_scan_code_l/_07_ ), .A2(\u_scan_code_l/_03_ ), .ZN(\u_scan_code_l/_08_ ) );
INV_X16 \u_scan_code_l/_47_ ( .A(\u_scan_code_l/_03_ ), .ZN(\u_scan_code_l/_09_ ) );
NOR2_X2 \u_scan_code_l/_48_ ( .A1(\u_scan_code_l/_09_ ), .A2(\u_scan_code_l/_02_ ), .ZN(\u_scan_code_l/_10_ ) );
OR3_X4 \u_scan_code_l/_49_ ( .A1(\u_scan_code_l/_06_ ), .A2(\u_scan_code_l/_08_ ), .A3(\u_scan_code_l/_10_ ), .ZN(\u_scan_code_l/_11_ ) );
INV_X32 \u_scan_code_l/_50_ ( .A(\u_scan_code_l/_00_ ), .ZN(\u_scan_code_l/_12_ ) );
NOR2_X2 \u_scan_code_l/_51_ ( .A1(\u_scan_code_l/_12_ ), .A2(\u_scan_code_l/_01_ ), .ZN(\u_scan_code_l/_13_ ) );
NOR2_X4 \u_scan_code_l/_52_ ( .A1(\u_scan_code_l/_03_ ), .A2(\u_scan_code_l/_02_ ), .ZN(\u_scan_code_l/_14_ ) );
AND2_X1 \u_scan_code_l/_53_ ( .A1(\u_scan_code_l/_13_ ), .A2(\u_scan_code_l/_14_ ), .ZN(\u_scan_code_l/_15_ ) );
INV_X1 \u_scan_code_l/_54_ ( .A(\u_scan_code_l/_15_ ), .ZN(\u_scan_code_l/_16_ ) );
INV_X1 \u_scan_code_l/_55_ ( .A(\u_scan_code_l/_04_ ), .ZN(\u_scan_code_l/_17_ ) );
AND2_X4 \u_scan_code_l/_56_ ( .A1(\u_scan_code_l/_01_ ), .A2(\u_scan_code_l/_00_ ), .ZN(\u_scan_code_l/_18_ ) );
AOI21_X1 \u_scan_code_l/_57_ ( .A(\u_scan_code_l/_17_ ), .B1(\u_scan_code_l/_08_ ), .B2(\u_scan_code_l/_18_ ), .ZN(\u_scan_code_l/_19_ ) );
NAND3_X1 \u_scan_code_l/_58_ ( .A1(\u_scan_code_l/_11_ ), .A2(\u_scan_code_l/_16_ ), .A3(\u_scan_code_l/_19_ ), .ZN(\u_scan_code_l/_35_ ) );
NAND2_X1 \u_scan_code_l/_59_ ( .A1(\u_scan_code_l/_06_ ), .A2(\u_scan_code_l/_14_ ), .ZN(\u_scan_code_l/_20_ ) );
AND2_X2 \u_scan_code_l/_60_ ( .A1(\u_scan_code_l/_03_ ), .A2(\u_scan_code_l/_02_ ), .ZN(\u_scan_code_l/_21_ ) );
NAND2_X1 \u_scan_code_l/_61_ ( .A1(\u_scan_code_l/_13_ ), .A2(\u_scan_code_l/_21_ ), .ZN(\u_scan_code_l/_22_ ) );
NAND3_X1 \u_scan_code_l/_62_ ( .A1(\u_scan_code_l/_19_ ), .A2(\u_scan_code_l/_20_ ), .A3(\u_scan_code_l/_22_ ), .ZN(\u_scan_code_l/_36_ ) );
NOR3_X1 \u_scan_code_l/_63_ ( .A1(\u_scan_code_l/_07_ ), .A2(\u_scan_code_l/_03_ ), .A3(\u_scan_code_l/_01_ ), .ZN(\u_scan_code_l/_23_ ) );
AOI21_X1 \u_scan_code_l/_64_ ( .A(\u_scan_code_l/_23_ ), .B1(\u_scan_code_l/_08_ ), .B2(\u_scan_code_l/_18_ ), .ZN(\u_scan_code_l/_24_ ) );
NAND3_X1 \u_scan_code_l/_65_ ( .A1(\u_scan_code_l/_09_ ), .A2(\u_scan_code_l/_07_ ), .A3(\u_scan_code_l/_00_ ), .ZN(\u_scan_code_l/_25_ ) );
NAND2_X1 \u_scan_code_l/_66_ ( .A1(\u_scan_code_l/_13_ ), .A2(\u_scan_code_l/_10_ ), .ZN(\u_scan_code_l/_26_ ) );
NAND4_X1 \u_scan_code_l/_67_ ( .A1(\u_scan_code_l/_24_ ), .A2(\u_scan_code_l/_04_ ), .A3(\u_scan_code_l/_25_ ), .A4(\u_scan_code_l/_26_ ), .ZN(\u_scan_code_l/_37_ ) );
NAND3_X1 \u_scan_code_l/_68_ ( .A1(\u_scan_code_l/_10_ ), .A2(\u_scan_code_l/_01_ ), .A3(\u_scan_code_l/_12_ ), .ZN(\u_scan_code_l/_27_ ) );
AOI22_X1 \u_scan_code_l/_69_ ( .A1(\u_scan_code_l/_08_ ), .A2(\u_scan_code_l/_05_ ), .B1(\u_scan_code_l/_18_ ), .B2(\u_scan_code_l/_21_ ), .ZN(\u_scan_code_l/_28_ ) );
NAND4_X1 \u_scan_code_l/_70_ ( .A1(\u_scan_code_l/_16_ ), .A2(\u_scan_code_l/_19_ ), .A3(\u_scan_code_l/_27_ ), .A4(\u_scan_code_l/_28_ ), .ZN(\u_scan_code_l/_38_ ) );
OAI21_X1 \u_scan_code_l/_71_ ( .A(\u_scan_code_l/_21_ ), .B1(\u_scan_code_l/_01_ ), .B2(\u_scan_code_l/_12_ ), .ZN(\u_scan_code_l/_29_ ) );
NAND3_X1 \u_scan_code_l/_72_ ( .A1(\u_scan_code_l/_14_ ), .A2(\u_scan_code_l/_01_ ), .A3(\u_scan_code_l/_12_ ), .ZN(\u_scan_code_l/_30_ ) );
NAND3_X1 \u_scan_code_l/_73_ ( .A1(\u_scan_code_l/_29_ ), .A2(\u_scan_code_l/_30_ ), .A3(\u_scan_code_l/_04_ ), .ZN(\u_scan_code_l/_39_ ) );
AND2_X1 \u_scan_code_l/_74_ ( .A1(\u_scan_code_l/_12_ ), .A2(\u_scan_code_l/_01_ ), .ZN(\u_scan_code_l/_31_ ) );
OAI21_X1 \u_scan_code_l/_75_ ( .A(\u_scan_code_l/_08_ ), .B1(\u_scan_code_l/_31_ ), .B2(\u_scan_code_l/_13_ ), .ZN(\u_scan_code_l/_32_ ) );
NAND2_X1 \u_scan_code_l/_76_ ( .A1(\u_scan_code_l/_10_ ), .A2(\u_scan_code_l/_18_ ), .ZN(\u_scan_code_l/_33_ ) );
NAND4_X1 \u_scan_code_l/_77_ ( .A1(\u_scan_code_l/_32_ ), .A2(\u_scan_code_l/_04_ ), .A3(\u_scan_code_l/_29_ ), .A4(\u_scan_code_l/_33_ ), .ZN(\u_scan_code_l/_40_ ) );
AOI22_X1 \u_scan_code_l/_78_ ( .A1(\u_scan_code_l/_14_ ), .A2(\u_scan_code_l/_13_ ), .B1(\u_scan_code_l/_08_ ), .B2(\u_scan_code_l/_05_ ), .ZN(\u_scan_code_l/_34_ ) );
NAND4_X1 \u_scan_code_l/_79_ ( .A1(\u_scan_code_l/_34_ ), .A2(\u_scan_code_l/_04_ ), .A3(\u_scan_code_l/_22_ ), .A4(\u_scan_code_l/_33_ ), .ZN(\u_scan_code_l/_41_ ) );
LOGIC1_X1 \u_scan_code_l/_80_ ( .Z(\u_scan_code_l/_42_ ) );
BUF_X1 \u_scan_code_l/_81_ ( .A(\u_scan_code_l/_42_ ), .Z(\scan_code_seg [0] ) );
BUF_X1 \u_scan_code_l/_82_ ( .A(\scan_code_buf [3] ), .Z(\u_scan_code_l/_03_ ) );
BUF_X1 \u_scan_code_l/_83_ ( .A(\scan_code_buf [2] ), .Z(\u_scan_code_l/_02_ ) );
BUF_X1 \u_scan_code_l/_84_ ( .A(\scan_code_buf [1] ), .Z(\u_scan_code_l/_01_ ) );
BUF_X1 \u_scan_code_l/_85_ ( .A(\scan_code_buf [0] ), .Z(\u_scan_code_l/_00_ ) );
BUF_X1 \u_scan_code_l/_86_ ( .A(display_en ), .Z(\u_scan_code_l/_04_ ) );
BUF_X1 \u_scan_code_l/_87_ ( .A(\u_scan_code_l/_35_ ), .Z(\scan_code_seg [1] ) );
BUF_X1 \u_scan_code_l/_88_ ( .A(\u_scan_code_l/_36_ ), .Z(\scan_code_seg [2] ) );
BUF_X1 \u_scan_code_l/_89_ ( .A(\u_scan_code_l/_37_ ), .Z(\scan_code_seg [3] ) );
BUF_X1 \u_scan_code_l/_90_ ( .A(\u_scan_code_l/_38_ ), .Z(\scan_code_seg [4] ) );
BUF_X1 \u_scan_code_l/_91_ ( .A(\u_scan_code_l/_39_ ), .Z(\scan_code_seg [5] ) );
BUF_X1 \u_scan_code_l/_92_ ( .A(\u_scan_code_l/_40_ ), .Z(\scan_code_seg [6] ) );
BUF_X1 \u_scan_code_l/_93_ ( .A(\u_scan_code_l/_41_ ), .Z(\scan_code_seg [7] ) );

endmodule
