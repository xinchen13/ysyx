module bitrev (
    input  sck,
    input  ss,
    input  mosi,
    output miso
);


    endmodule
