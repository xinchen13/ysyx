//Generate the verilog at 2024-07-13T10:15:50
module top (
clk,
rst_n,
data,
segment_dis
);

input clk ;
input rst_n ;
input [7:0] data ;
output [15:0] segment_dis ;

wire \u_lfsr/_00_ ;
wire \u_lfsr/_01_ ;
wire \u_lfsr/_02_ ;
wire \u_lfsr/_03_ ;
wire \u_lfsr/_04_ ;
wire \u_lfsr/_05_ ;
wire \u_lfsr/_06_ ;
wire \u_lfsr/_07_ ;
wire \u_lfsr/_08_ ;
wire \u_lfsr/_09_ ;
wire \u_lfsr/_10_ ;
wire \u_lfsr/_11_ ;
wire \u_lfsr/_12_ ;
wire \u_lfsr/_13_ ;
wire \u_lfsr/_14_ ;
wire \u_lfsr/_15_ ;
wire \u_lfsr/_16_ ;
wire \u_lfsr/_17_ ;
wire \u_lfsr/_18_ ;
wire \u_lfsr/_19_ ;
wire \u_lfsr/_20_ ;
wire \u_lfsr/_21_ ;
wire \u_lfsr/_22_ ;
wire \u_lfsr/_23_ ;
wire \u_lfsr/_24_ ;
wire \u_lfsr/_25_ ;
wire \u_lfsr/_26_ ;
wire \u_lfsr/_27_ ;
wire \u_lfsr/_28_ ;
wire \u_lfsr/_29_ ;
wire \u_lfsr/_30_ ;
wire \u_lfsr/_31_ ;
wire \u_lfsr/_32_ ;
wire \u_lfsr/_33_ ;
wire \u_lfsr/_34_ ;
wire \u_lfsr/_35_ ;
wire \u_lfsr/_36_ ;
wire \u_lfsr/_37_ ;
wire \u_lfsr/_38_ ;
wire \u_lfsr/_39_ ;
wire \u_lfsr/_40_ ;
wire \u_lfsr/_41_ ;
wire \u_lfsr/_42_ ;
wire \u_lfsr/_43_ ;
wire \u_seg1/_00_ ;
wire \u_seg1/_01_ ;
wire \u_seg1/_02_ ;
wire \u_seg1/_03_ ;
wire \u_seg1/_04_ ;
wire \u_seg1/_05_ ;
wire \u_seg1/_06_ ;
wire \u_seg1/_07_ ;
wire \u_seg1/_08_ ;
wire \u_seg1/_09_ ;
wire \u_seg1/_10_ ;
wire \u_seg1/_11_ ;
wire \u_seg1/_12_ ;
wire \u_seg1/_13_ ;
wire \u_seg1/_14_ ;
wire \u_seg1/_15_ ;
wire \u_seg1/_16_ ;
wire \u_seg1/_17_ ;
wire \u_seg1/_18_ ;
wire \u_seg1/_19_ ;
wire \u_seg1/_20_ ;
wire \u_seg1/_21_ ;
wire \u_seg1/_22_ ;
wire \u_seg1/_23_ ;
wire \u_seg1/_24_ ;
wire \u_seg1/_25_ ;
wire \u_seg1/_26_ ;
wire \u_seg1/_27_ ;
wire \u_seg1/_28_ ;
wire \u_seg1/_29_ ;
wire \u_seg1/_30_ ;
wire \u_seg1/_31_ ;
wire \u_seg1/_32_ ;
wire \u_seg1/_33_ ;
wire \u_seg1/_34_ ;
wire \u_seg1/_35_ ;
wire \u_seg1/_36_ ;
wire \u_seg1/_37_ ;
wire \u_seg1/_38_ ;
wire \u_seg2/_00_ ;
wire \u_seg2/_01_ ;
wire \u_seg2/_02_ ;
wire \u_seg2/_03_ ;
wire \u_seg2/_04_ ;
wire \u_seg2/_05_ ;
wire \u_seg2/_06_ ;
wire \u_seg2/_07_ ;
wire \u_seg2/_08_ ;
wire \u_seg2/_09_ ;
wire \u_seg2/_10_ ;
wire \u_seg2/_11_ ;
wire \u_seg2/_12_ ;
wire \u_seg2/_13_ ;
wire \u_seg2/_14_ ;
wire \u_seg2/_15_ ;
wire \u_seg2/_16_ ;
wire \u_seg2/_17_ ;
wire \u_seg2/_18_ ;
wire \u_seg2/_19_ ;
wire \u_seg2/_20_ ;
wire \u_seg2/_21_ ;
wire \u_seg2/_22_ ;
wire \u_seg2/_23_ ;
wire \u_seg2/_24_ ;
wire \u_seg2/_25_ ;
wire \u_seg2/_26_ ;
wire \u_seg2/_27_ ;
wire \u_seg2/_28_ ;
wire \u_seg2/_29_ ;
wire \u_seg2/_30_ ;
wire \u_seg2/_31_ ;
wire \u_seg2/_32_ ;
wire \u_seg2/_33_ ;
wire \u_seg2/_34_ ;
wire \u_seg2/_35_ ;
wire \u_seg2/_36_ ;
wire \u_seg2/_37_ ;
wire \u_seg2/_38_ ;
wire rst_n ;
wire clk ;
wire \bcd[0] ;
wire \bcd[1] ;
wire \bcd[2] ;
wire \bcd[3] ;
wire \bcd[4] ;
wire \bcd[5] ;
wire \bcd[6] ;
wire \bcd[7] ;
wire \data[0] ;
wire \data[1] ;
wire \data[2] ;
wire \data[3] ;
wire \data[4] ;
wire \data[5] ;
wire \data[6] ;
wire \data[7] ;
wire \segment_dis[0] ;
wire \segment_dis[1] ;
wire \segment_dis[2] ;
wire \segment_dis[3] ;
wire \segment_dis[4] ;
wire \segment_dis[5] ;
wire \segment_dis[6] ;
wire \segment_dis[7] ;
wire \segment_dis[8] ;
wire \segment_dis[9] ;
wire \segment_dis[10] ;
wire \segment_dis[11] ;
wire \segment_dis[12] ;
wire \segment_dis[13] ;
wire \segment_dis[14] ;
wire \segment_dis[15] ;

assign \data[0] = data[0] ;
assign \data[1] = data[1] ;
assign \data[2] = data[2] ;
assign \data[3] = data[3] ;
assign \data[4] = data[4] ;
assign \data[5] = data[5] ;
assign \data[6] = data[6] ;
assign \data[7] = data[7] ;
assign segment_dis[0] = \segment_dis[0] ;
assign segment_dis[1] = \segment_dis[1] ;
assign segment_dis[2] = \segment_dis[2] ;
assign segment_dis[3] = \segment_dis[3] ;
assign segment_dis[4] = \segment_dis[4] ;
assign segment_dis[5] = \segment_dis[5] ;
assign segment_dis[6] = \segment_dis[6] ;
assign segment_dis[7] = \segment_dis[7] ;
assign segment_dis[8] = \segment_dis[8] ;
assign segment_dis[9] = \segment_dis[9] ;
assign segment_dis[10] = \segment_dis[10] ;
assign segment_dis[11] = \segment_dis[11] ;
assign segment_dis[12] = \segment_dis[12] ;
assign segment_dis[13] = \segment_dis[13] ;
assign segment_dis[14] = \segment_dis[14] ;
assign segment_dis[15] = \segment_dis[15] ;

MUX2_X1 \u_lfsr/_44_ ( .A(\u_lfsr/_16_ ), .B(\u_lfsr/_25_ ), .S(\u_lfsr/_35_ ), .Z(\u_lfsr/_08_ ) );
MUX2_X1 \u_lfsr/_45_ ( .A(\u_lfsr/_17_ ), .B(\u_lfsr/_26_ ), .S(\u_lfsr/_35_ ), .Z(\u_lfsr/_09_ ) );
MUX2_X1 \u_lfsr/_46_ ( .A(\u_lfsr/_18_ ), .B(\u_lfsr/_27_ ), .S(\u_lfsr/_35_ ), .Z(\u_lfsr/_10_ ) );
MUX2_X1 \u_lfsr/_47_ ( .A(\u_lfsr/_19_ ), .B(\u_lfsr/_28_ ), .S(\u_lfsr/_35_ ), .Z(\u_lfsr/_11_ ) );
MUX2_X1 \u_lfsr/_48_ ( .A(\u_lfsr/_20_ ), .B(\u_lfsr/_29_ ), .S(\u_lfsr/_35_ ), .Z(\u_lfsr/_12_ ) );
MUX2_X1 \u_lfsr/_49_ ( .A(\u_lfsr/_21_ ), .B(\u_lfsr/_30_ ), .S(\u_lfsr/_35_ ), .Z(\u_lfsr/_13_ ) );
MUX2_X1 \u_lfsr/_50_ ( .A(\u_lfsr/_22_ ), .B(\u_lfsr/_31_ ), .S(\u_lfsr/_35_ ), .Z(\u_lfsr/_14_ ) );
XOR2_X2 \u_lfsr/_51_ ( .A(\u_lfsr/_28_ ), .B(\u_lfsr/_24_ ), .Z(\u_lfsr/_32_ ) );
XNOR2_X2 \u_lfsr/_52_ ( .A(\u_lfsr/_26_ ), .B(\u_lfsr/_27_ ), .ZN(\u_lfsr/_33_ ) );
XNOR2_X1 \u_lfsr/_53_ ( .A(\u_lfsr/_32_ ), .B(\u_lfsr/_33_ ), .ZN(\u_lfsr/_34_ ) );
MUX2_X2 \u_lfsr/_54_ ( .A(\u_lfsr/_23_ ), .B(\u_lfsr/_34_ ), .S(\u_lfsr/_35_ ), .Z(\u_lfsr/_15_ ) );
BUF_X1 \u_lfsr/_55_ ( .A(\data[0] ), .Z(\u_lfsr/_16_ ) );
BUF_X1 \u_lfsr/_56_ ( .A(\bcd[1] ), .Z(\u_lfsr/_25_ ) );
BUF_X1 \u_lfsr/_57_ ( .A(rst_n ), .Z(\u_lfsr/_35_ ) );
BUF_X1 \u_lfsr/_58_ ( .A(\u_lfsr/_08_ ), .Z(\u_lfsr/_00_ ) );
BUF_X1 \u_lfsr/_59_ ( .A(\data[1] ), .Z(\u_lfsr/_17_ ) );
BUF_X1 \u_lfsr/_60_ ( .A(\bcd[2] ), .Z(\u_lfsr/_26_ ) );
BUF_X1 \u_lfsr/_61_ ( .A(\u_lfsr/_09_ ), .Z(\u_lfsr/_01_ ) );
BUF_X1 \u_lfsr/_62_ ( .A(\data[2] ), .Z(\u_lfsr/_18_ ) );
BUF_X1 \u_lfsr/_63_ ( .A(\bcd[3] ), .Z(\u_lfsr/_27_ ) );
BUF_X1 \u_lfsr/_64_ ( .A(\u_lfsr/_10_ ), .Z(\u_lfsr/_02_ ) );
BUF_X1 \u_lfsr/_65_ ( .A(\data[3] ), .Z(\u_lfsr/_19_ ) );
BUF_X1 \u_lfsr/_66_ ( .A(\bcd[4] ), .Z(\u_lfsr/_28_ ) );
BUF_X1 \u_lfsr/_67_ ( .A(\u_lfsr/_11_ ), .Z(\u_lfsr/_03_ ) );
BUF_X1 \u_lfsr/_68_ ( .A(\data[4] ), .Z(\u_lfsr/_20_ ) );
BUF_X1 \u_lfsr/_69_ ( .A(\bcd[5] ), .Z(\u_lfsr/_29_ ) );
BUF_X1 \u_lfsr/_70_ ( .A(\u_lfsr/_12_ ), .Z(\u_lfsr/_04_ ) );
BUF_X1 \u_lfsr/_71_ ( .A(\data[5] ), .Z(\u_lfsr/_21_ ) );
BUF_X1 \u_lfsr/_72_ ( .A(\bcd[6] ), .Z(\u_lfsr/_30_ ) );
BUF_X1 \u_lfsr/_73_ ( .A(\u_lfsr/_13_ ), .Z(\u_lfsr/_05_ ) );
BUF_X1 \u_lfsr/_74_ ( .A(\data[6] ), .Z(\u_lfsr/_22_ ) );
BUF_X1 \u_lfsr/_75_ ( .A(\bcd[7] ), .Z(\u_lfsr/_31_ ) );
BUF_X1 \u_lfsr/_76_ ( .A(\u_lfsr/_14_ ), .Z(\u_lfsr/_06_ ) );
BUF_X1 \u_lfsr/_77_ ( .A(\bcd[0] ), .Z(\u_lfsr/_24_ ) );
BUF_X1 \u_lfsr/_78_ ( .A(\data[7] ), .Z(\u_lfsr/_23_ ) );
BUF_X1 \u_lfsr/_79_ ( .A(\u_lfsr/_15_ ), .Z(\u_lfsr/_07_ ) );
DFF_X1 \u_lfsr/_80_ ( .D(\u_lfsr/_00_ ), .CK(clk ), .Q(\bcd[0] ), .QN(\u_lfsr/_36_ ) );
DFF_X1 \u_lfsr/_81_ ( .D(\u_lfsr/_01_ ), .CK(clk ), .Q(\bcd[1] ), .QN(\u_lfsr/_37_ ) );
DFF_X1 \u_lfsr/_82_ ( .D(\u_lfsr/_02_ ), .CK(clk ), .Q(\bcd[2] ), .QN(\u_lfsr/_38_ ) );
DFF_X1 \u_lfsr/_83_ ( .D(\u_lfsr/_03_ ), .CK(clk ), .Q(\bcd[3] ), .QN(\u_lfsr/_39_ ) );
DFF_X1 \u_lfsr/_84_ ( .D(\u_lfsr/_04_ ), .CK(clk ), .Q(\bcd[4] ), .QN(\u_lfsr/_40_ ) );
DFF_X1 \u_lfsr/_85_ ( .D(\u_lfsr/_05_ ), .CK(clk ), .Q(\bcd[5] ), .QN(\u_lfsr/_41_ ) );
DFF_X1 \u_lfsr/_86_ ( .D(\u_lfsr/_06_ ), .CK(clk ), .Q(\bcd[6] ), .QN(\u_lfsr/_42_ ) );
DFF_X1 \u_lfsr/_87_ ( .D(\u_lfsr/_07_ ), .CK(clk ), .Q(\bcd[7] ), .QN(\u_lfsr/_43_ ) );
INV_X16 \u_seg1/_39_ ( .A(\u_seg1/_02_ ), .ZN(\u_seg1/_04_ ) );
NOR2_X4 \u_seg1/_40_ ( .A1(\u_seg1/_04_ ), .A2(\u_seg1/_03_ ), .ZN(\u_seg1/_05_ ) );
AND2_X4 \u_seg1/_41_ ( .A1(\u_seg1/_01_ ), .A2(\u_seg1/_00_ ), .ZN(\u_seg1/_06_ ) );
AND2_X4 \u_seg1/_42_ ( .A1(\u_seg1/_05_ ), .A2(\u_seg1/_06_ ), .ZN(\u_seg1/_07_ ) );
NOR2_X4 \u_seg1/_43_ ( .A1(\u_seg1/_03_ ), .A2(\u_seg1/_02_ ), .ZN(\u_seg1/_08_ ) );
INV_X16 \u_seg1/_44_ ( .A(\u_seg1/_00_ ), .ZN(\u_seg1/_09_ ) );
NOR2_X2 \u_seg1/_45_ ( .A1(\u_seg1/_09_ ), .A2(\u_seg1/_01_ ), .ZN(\u_seg1/_10_ ) );
AOI21_X4 \u_seg1/_46_ ( .A(\u_seg1/_07_ ), .B1(\u_seg1/_08_ ), .B2(\u_seg1/_10_ ), .ZN(\u_seg1/_11_ ) );
INV_X1 \u_seg1/_47_ ( .A(\u_seg1/_05_ ), .ZN(\u_seg1/_12_ ) );
INV_X1 \u_seg1/_48_ ( .A(\u_seg1/_03_ ), .ZN(\u_seg1/_13_ ) );
NOR2_X1 \u_seg1/_49_ ( .A1(\u_seg1/_13_ ), .A2(\u_seg1/_02_ ), .ZN(\u_seg1/_14_ ) );
INV_X1 \u_seg1/_50_ ( .A(\u_seg1/_14_ ), .ZN(\u_seg1/_15_ ) );
NOR2_X1 \u_seg1/_51_ ( .A1(\u_seg1/_01_ ), .A2(\u_seg1/_00_ ), .ZN(\u_seg1/_16_ ) );
NAND3_X1 \u_seg1/_52_ ( .A1(\u_seg1/_12_ ), .A2(\u_seg1/_15_ ), .A3(\u_seg1/_16_ ), .ZN(\u_seg1/_17_ ) );
NAND2_X1 \u_seg1/_53_ ( .A1(\u_seg1/_11_ ), .A2(\u_seg1/_17_ ), .ZN(\u_seg1/_31_ ) );
AND2_X2 \u_seg1/_54_ ( .A1(\u_seg1/_03_ ), .A2(\u_seg1/_02_ ), .ZN(\u_seg1/_18_ ) );
NAND2_X1 \u_seg1/_55_ ( .A1(\u_seg1/_10_ ), .A2(\u_seg1/_18_ ), .ZN(\u_seg1/_19_ ) );
INV_X1 \u_seg1/_56_ ( .A(\u_seg1/_08_ ), .ZN(\u_seg1/_20_ ) );
INV_X1 \u_seg1/_57_ ( .A(\u_seg1/_06_ ), .ZN(\u_seg1/_21_ ) );
OAI221_X1 \u_seg1/_58_ ( .A(\u_seg1/_19_ ), .B1(\u_seg1/_20_ ), .B2(\u_seg1/_16_ ), .C1(\u_seg1/_12_ ), .C2(\u_seg1/_21_ ), .ZN(\u_seg1/_32_ ) );
INV_X32 \u_seg1/_59_ ( .A(\u_seg1/_01_ ), .ZN(\u_seg1/_22_ ) );
OAI211_X2 \u_seg1/_60_ ( .A(\u_seg1/_13_ ), .B(\u_seg1/_02_ ), .C1(\u_seg1/_22_ ), .C2(\u_seg1/_00_ ), .ZN(\u_seg1/_23_ ) );
NAND4_X1 \u_seg1/_61_ ( .A1(\u_seg1/_04_ ), .A2(\u_seg1/_22_ ), .A3(\u_seg1/_03_ ), .A4(\u_seg1/_00_ ), .ZN(\u_seg1/_24_ ) );
OAI211_X2 \u_seg1/_62_ ( .A(\u_seg1/_23_ ), .B(\u_seg1/_24_ ), .C1(\u_seg1/_20_ ), .C2(\u_seg1/_09_ ), .ZN(\u_seg1/_33_ ) );
AOI22_X1 \u_seg1/_63_ ( .A1(\u_seg1/_05_ ), .A2(\u_seg1/_16_ ), .B1(\u_seg1/_06_ ), .B2(\u_seg1/_18_ ), .ZN(\u_seg1/_25_ ) );
NOR2_X1 \u_seg1/_64_ ( .A1(\u_seg1/_22_ ), .A2(\u_seg1/_00_ ), .ZN(\u_seg1/_26_ ) );
INV_X1 \u_seg1/_65_ ( .A(\u_seg1/_26_ ), .ZN(\u_seg1/_27_ ) );
OAI211_X2 \u_seg1/_66_ ( .A(\u_seg1/_11_ ), .B(\u_seg1/_25_ ), .C1(\u_seg1/_15_ ), .C2(\u_seg1/_27_ ), .ZN(\u_seg1/_34_ ) );
OAI21_X1 \u_seg1/_67_ ( .A(\u_seg1/_18_ ), .B1(\u_seg1/_01_ ), .B2(\u_seg1/_09_ ), .ZN(\u_seg1/_28_ ) );
OAI21_X1 \u_seg1/_68_ ( .A(\u_seg1/_28_ ), .B1(\u_seg1/_27_ ), .B2(\u_seg1/_20_ ), .ZN(\u_seg1/_35_ ) );
OAI21_X1 \u_seg1/_69_ ( .A(\u_seg1/_05_ ), .B1(\u_seg1/_10_ ), .B2(\u_seg1/_26_ ), .ZN(\u_seg1/_29_ ) );
OAI211_X2 \u_seg1/_70_ ( .A(\u_seg1/_29_ ), .B(\u_seg1/_28_ ), .C1(\u_seg1/_21_ ), .C2(\u_seg1/_15_ ), .ZN(\u_seg1/_36_ ) );
AOI22_X1 \u_seg1/_71_ ( .A1(\u_seg1/_08_ ), .A2(\u_seg1/_10_ ), .B1(\u_seg1/_05_ ), .B2(\u_seg1/_16_ ), .ZN(\u_seg1/_30_ ) );
OAI211_X2 \u_seg1/_72_ ( .A(\u_seg1/_30_ ), .B(\u_seg1/_19_ ), .C1(\u_seg1/_21_ ), .C2(\u_seg1/_15_ ), .ZN(\u_seg1/_37_ ) );
LOGIC1_X1 \u_seg1/_73_ ( .Z(\u_seg1/_38_ ) );
BUF_X1 \u_seg1/_74_ ( .A(\u_seg1/_38_ ), .Z(\segment_dis[0] ) );
BUF_X1 \u_seg1/_75_ ( .A(\bcd[3] ), .Z(\u_seg1/_03_ ) );
BUF_X1 \u_seg1/_76_ ( .A(\bcd[2] ), .Z(\u_seg1/_02_ ) );
BUF_X1 \u_seg1/_77_ ( .A(\bcd[1] ), .Z(\u_seg1/_01_ ) );
BUF_X1 \u_seg1/_78_ ( .A(\bcd[0] ), .Z(\u_seg1/_00_ ) );
BUF_X1 \u_seg1/_79_ ( .A(\u_seg1/_31_ ), .Z(\segment_dis[1] ) );
BUF_X1 \u_seg1/_80_ ( .A(\u_seg1/_32_ ), .Z(\segment_dis[2] ) );
BUF_X1 \u_seg1/_81_ ( .A(\u_seg1/_33_ ), .Z(\segment_dis[3] ) );
BUF_X1 \u_seg1/_82_ ( .A(\u_seg1/_34_ ), .Z(\segment_dis[4] ) );
BUF_X1 \u_seg1/_83_ ( .A(\u_seg1/_35_ ), .Z(\segment_dis[5] ) );
BUF_X1 \u_seg1/_84_ ( .A(\u_seg1/_36_ ), .Z(\segment_dis[6] ) );
BUF_X1 \u_seg1/_85_ ( .A(\u_seg1/_37_ ), .Z(\segment_dis[7] ) );
INV_X16 \u_seg2/_39_ ( .A(\u_seg2/_02_ ), .ZN(\u_seg2/_04_ ) );
NOR2_X4 \u_seg2/_40_ ( .A1(\u_seg2/_04_ ), .A2(\u_seg2/_03_ ), .ZN(\u_seg2/_05_ ) );
AND2_X4 \u_seg2/_41_ ( .A1(\u_seg2/_01_ ), .A2(\u_seg2/_00_ ), .ZN(\u_seg2/_06_ ) );
AND2_X4 \u_seg2/_42_ ( .A1(\u_seg2/_05_ ), .A2(\u_seg2/_06_ ), .ZN(\u_seg2/_07_ ) );
NOR2_X4 \u_seg2/_43_ ( .A1(\u_seg2/_03_ ), .A2(\u_seg2/_02_ ), .ZN(\u_seg2/_08_ ) );
INV_X16 \u_seg2/_44_ ( .A(\u_seg2/_00_ ), .ZN(\u_seg2/_09_ ) );
NOR2_X2 \u_seg2/_45_ ( .A1(\u_seg2/_09_ ), .A2(\u_seg2/_01_ ), .ZN(\u_seg2/_10_ ) );
AOI21_X4 \u_seg2/_46_ ( .A(\u_seg2/_07_ ), .B1(\u_seg2/_08_ ), .B2(\u_seg2/_10_ ), .ZN(\u_seg2/_11_ ) );
INV_X1 \u_seg2/_47_ ( .A(\u_seg2/_05_ ), .ZN(\u_seg2/_12_ ) );
INV_X1 \u_seg2/_48_ ( .A(\u_seg2/_03_ ), .ZN(\u_seg2/_13_ ) );
NOR2_X1 \u_seg2/_49_ ( .A1(\u_seg2/_13_ ), .A2(\u_seg2/_02_ ), .ZN(\u_seg2/_14_ ) );
INV_X1 \u_seg2/_50_ ( .A(\u_seg2/_14_ ), .ZN(\u_seg2/_15_ ) );
NOR2_X1 \u_seg2/_51_ ( .A1(\u_seg2/_01_ ), .A2(\u_seg2/_00_ ), .ZN(\u_seg2/_16_ ) );
NAND3_X1 \u_seg2/_52_ ( .A1(\u_seg2/_12_ ), .A2(\u_seg2/_15_ ), .A3(\u_seg2/_16_ ), .ZN(\u_seg2/_17_ ) );
NAND2_X1 \u_seg2/_53_ ( .A1(\u_seg2/_11_ ), .A2(\u_seg2/_17_ ), .ZN(\u_seg2/_31_ ) );
AND2_X2 \u_seg2/_54_ ( .A1(\u_seg2/_03_ ), .A2(\u_seg2/_02_ ), .ZN(\u_seg2/_18_ ) );
NAND2_X1 \u_seg2/_55_ ( .A1(\u_seg2/_10_ ), .A2(\u_seg2/_18_ ), .ZN(\u_seg2/_19_ ) );
INV_X1 \u_seg2/_56_ ( .A(\u_seg2/_08_ ), .ZN(\u_seg2/_20_ ) );
INV_X1 \u_seg2/_57_ ( .A(\u_seg2/_06_ ), .ZN(\u_seg2/_21_ ) );
OAI221_X1 \u_seg2/_58_ ( .A(\u_seg2/_19_ ), .B1(\u_seg2/_20_ ), .B2(\u_seg2/_16_ ), .C1(\u_seg2/_12_ ), .C2(\u_seg2/_21_ ), .ZN(\u_seg2/_32_ ) );
INV_X32 \u_seg2/_59_ ( .A(\u_seg2/_01_ ), .ZN(\u_seg2/_22_ ) );
OAI211_X2 \u_seg2/_60_ ( .A(\u_seg2/_13_ ), .B(\u_seg2/_02_ ), .C1(\u_seg2/_22_ ), .C2(\u_seg2/_00_ ), .ZN(\u_seg2/_23_ ) );
NAND4_X1 \u_seg2/_61_ ( .A1(\u_seg2/_04_ ), .A2(\u_seg2/_22_ ), .A3(\u_seg2/_03_ ), .A4(\u_seg2/_00_ ), .ZN(\u_seg2/_24_ ) );
OAI211_X2 \u_seg2/_62_ ( .A(\u_seg2/_23_ ), .B(\u_seg2/_24_ ), .C1(\u_seg2/_20_ ), .C2(\u_seg2/_09_ ), .ZN(\u_seg2/_33_ ) );
AOI22_X1 \u_seg2/_63_ ( .A1(\u_seg2/_05_ ), .A2(\u_seg2/_16_ ), .B1(\u_seg2/_06_ ), .B2(\u_seg2/_18_ ), .ZN(\u_seg2/_25_ ) );
NOR2_X1 \u_seg2/_64_ ( .A1(\u_seg2/_22_ ), .A2(\u_seg2/_00_ ), .ZN(\u_seg2/_26_ ) );
INV_X1 \u_seg2/_65_ ( .A(\u_seg2/_26_ ), .ZN(\u_seg2/_27_ ) );
OAI211_X2 \u_seg2/_66_ ( .A(\u_seg2/_11_ ), .B(\u_seg2/_25_ ), .C1(\u_seg2/_15_ ), .C2(\u_seg2/_27_ ), .ZN(\u_seg2/_34_ ) );
OAI21_X1 \u_seg2/_67_ ( .A(\u_seg2/_18_ ), .B1(\u_seg2/_01_ ), .B2(\u_seg2/_09_ ), .ZN(\u_seg2/_28_ ) );
OAI21_X1 \u_seg2/_68_ ( .A(\u_seg2/_28_ ), .B1(\u_seg2/_27_ ), .B2(\u_seg2/_20_ ), .ZN(\u_seg2/_35_ ) );
OAI21_X1 \u_seg2/_69_ ( .A(\u_seg2/_05_ ), .B1(\u_seg2/_10_ ), .B2(\u_seg2/_26_ ), .ZN(\u_seg2/_29_ ) );
OAI211_X2 \u_seg2/_70_ ( .A(\u_seg2/_29_ ), .B(\u_seg2/_28_ ), .C1(\u_seg2/_21_ ), .C2(\u_seg2/_15_ ), .ZN(\u_seg2/_36_ ) );
AOI22_X1 \u_seg2/_71_ ( .A1(\u_seg2/_08_ ), .A2(\u_seg2/_10_ ), .B1(\u_seg2/_05_ ), .B2(\u_seg2/_16_ ), .ZN(\u_seg2/_30_ ) );
OAI211_X2 \u_seg2/_72_ ( .A(\u_seg2/_30_ ), .B(\u_seg2/_19_ ), .C1(\u_seg2/_21_ ), .C2(\u_seg2/_15_ ), .ZN(\u_seg2/_37_ ) );
LOGIC1_X1 \u_seg2/_73_ ( .Z(\u_seg2/_38_ ) );
BUF_X1 \u_seg2/_74_ ( .A(\u_seg2/_38_ ), .Z(\segment_dis[8] ) );
BUF_X1 \u_seg2/_75_ ( .A(\bcd[7] ), .Z(\u_seg2/_03_ ) );
BUF_X1 \u_seg2/_76_ ( .A(\bcd[6] ), .Z(\u_seg2/_02_ ) );
BUF_X1 \u_seg2/_77_ ( .A(\bcd[5] ), .Z(\u_seg2/_01_ ) );
BUF_X1 \u_seg2/_78_ ( .A(\bcd[4] ), .Z(\u_seg2/_00_ ) );
BUF_X1 \u_seg2/_79_ ( .A(\u_seg2/_31_ ), .Z(\segment_dis[9] ) );
BUF_X1 \u_seg2/_80_ ( .A(\u_seg2/_32_ ), .Z(\segment_dis[10] ) );
BUF_X1 \u_seg2/_81_ ( .A(\u_seg2/_33_ ), .Z(\segment_dis[11] ) );
BUF_X1 \u_seg2/_82_ ( .A(\u_seg2/_34_ ), .Z(\segment_dis[12] ) );
BUF_X1 \u_seg2/_83_ ( .A(\u_seg2/_35_ ), .Z(\segment_dis[13] ) );
BUF_X1 \u_seg2/_84_ ( .A(\u_seg2/_36_ ), .Z(\segment_dis[14] ) );
BUF_X1 \u_seg2/_85_ ( .A(\u_seg2/_37_ ), .Z(\segment_dis[15] ) );

endmodule
