//Generate the verilog at 2024-08-23T20:33:42
module alu2 (
clk,
a,
b,
ctrl,
result
);

input clk ;
input [31:0] a ;
input [31:0] b ;
input [3:0] ctrl ;
output [31:0] result ;

wire _0000_ ;
wire _0001_ ;
wire _0002_ ;
wire _0003_ ;
wire _0004_ ;
wire _0005_ ;
wire _0006_ ;
wire _0007_ ;
wire _0008_ ;
wire _0009_ ;
wire _0010_ ;
wire _0011_ ;
wire _0012_ ;
wire _0013_ ;
wire _0014_ ;
wire _0015_ ;
wire _0016_ ;
wire _0017_ ;
wire _0018_ ;
wire _0019_ ;
wire _0020_ ;
wire _0021_ ;
wire _0022_ ;
wire _0023_ ;
wire _0024_ ;
wire _0025_ ;
wire _0026_ ;
wire _0027_ ;
wire _0028_ ;
wire _0029_ ;
wire _0030_ ;
wire _0031_ ;
wire _0032_ ;
wire _0033_ ;
wire _0034_ ;
wire _0035_ ;
wire _0036_ ;
wire _0037_ ;
wire _0038_ ;
wire _0039_ ;
wire _0040_ ;
wire _0041_ ;
wire _0042_ ;
wire _0043_ ;
wire _0044_ ;
wire _0045_ ;
wire _0046_ ;
wire _0047_ ;
wire _0048_ ;
wire _0049_ ;
wire _0050_ ;
wire _0051_ ;
wire _0052_ ;
wire _0053_ ;
wire _0054_ ;
wire _0055_ ;
wire _0056_ ;
wire _0057_ ;
wire _0058_ ;
wire _0059_ ;
wire _0060_ ;
wire _0061_ ;
wire _0062_ ;
wire _0063_ ;
wire _0064_ ;
wire _0065_ ;
wire _0066_ ;
wire _0067_ ;
wire _0068_ ;
wire _0069_ ;
wire _0070_ ;
wire _0071_ ;
wire _0072_ ;
wire _0073_ ;
wire _0074_ ;
wire _0075_ ;
wire _0076_ ;
wire _0077_ ;
wire _0078_ ;
wire _0079_ ;
wire _0080_ ;
wire _0081_ ;
wire _0082_ ;
wire _0083_ ;
wire _0084_ ;
wire _0085_ ;
wire _0086_ ;
wire _0087_ ;
wire _0088_ ;
wire _0089_ ;
wire _0090_ ;
wire _0091_ ;
wire _0092_ ;
wire _0093_ ;
wire _0094_ ;
wire _0095_ ;
wire _0096_ ;
wire _0097_ ;
wire _0098_ ;
wire _0099_ ;
wire _0100_ ;
wire _0101_ ;
wire _0102_ ;
wire _0103_ ;
wire _0104_ ;
wire _0105_ ;
wire _0106_ ;
wire _0107_ ;
wire _0108_ ;
wire _0109_ ;
wire _0110_ ;
wire _0111_ ;
wire _0112_ ;
wire _0113_ ;
wire _0114_ ;
wire _0115_ ;
wire _0116_ ;
wire _0117_ ;
wire _0118_ ;
wire _0119_ ;
wire _0120_ ;
wire _0121_ ;
wire _0122_ ;
wire _0123_ ;
wire _0124_ ;
wire _0125_ ;
wire _0126_ ;
wire _0127_ ;
wire _0128_ ;
wire _0129_ ;
wire _0130_ ;
wire _0131_ ;
wire _0132_ ;
wire _0133_ ;
wire _0134_ ;
wire _0135_ ;
wire _0136_ ;
wire _0137_ ;
wire _0138_ ;
wire _0139_ ;
wire _0140_ ;
wire _0141_ ;
wire _0142_ ;
wire _0143_ ;
wire _0144_ ;
wire _0145_ ;
wire _0146_ ;
wire _0147_ ;
wire _0148_ ;
wire _0149_ ;
wire _0150_ ;
wire _0151_ ;
wire _0152_ ;
wire _0153_ ;
wire _0154_ ;
wire _0155_ ;
wire _0156_ ;
wire _0157_ ;
wire _0158_ ;
wire _0159_ ;
wire _0160_ ;
wire _0161_ ;
wire _0162_ ;
wire _0163_ ;
wire _0164_ ;
wire _0165_ ;
wire _0166_ ;
wire _0167_ ;
wire _0168_ ;
wire _0169_ ;
wire _0170_ ;
wire _0171_ ;
wire _0172_ ;
wire _0173_ ;
wire _0174_ ;
wire _0175_ ;
wire _0176_ ;
wire _0177_ ;
wire _0178_ ;
wire _0179_ ;
wire _0180_ ;
wire _0181_ ;
wire _0182_ ;
wire _0183_ ;
wire _0184_ ;
wire _0185_ ;
wire _0186_ ;
wire _0187_ ;
wire _0188_ ;
wire _0189_ ;
wire _0190_ ;
wire _0191_ ;
wire _0192_ ;
wire _0193_ ;
wire _0194_ ;
wire _0195_ ;
wire _0196_ ;
wire _0197_ ;
wire _0198_ ;
wire _0199_ ;
wire _0200_ ;
wire _0201_ ;
wire _0202_ ;
wire _0203_ ;
wire _0204_ ;
wire _0205_ ;
wire _0206_ ;
wire _0207_ ;
wire _0208_ ;
wire _0209_ ;
wire _0210_ ;
wire _0211_ ;
wire _0212_ ;
wire _0213_ ;
wire _0214_ ;
wire _0215_ ;
wire _0216_ ;
wire _0217_ ;
wire _0218_ ;
wire _0219_ ;
wire _0220_ ;
wire _0221_ ;
wire _0222_ ;
wire _0223_ ;
wire _0224_ ;
wire _0225_ ;
wire _0226_ ;
wire _0227_ ;
wire _0228_ ;
wire _0229_ ;
wire _0230_ ;
wire _0231_ ;
wire _0232_ ;
wire _0233_ ;
wire _0234_ ;
wire _0235_ ;
wire _0236_ ;
wire _0237_ ;
wire _0238_ ;
wire _0239_ ;
wire _0240_ ;
wire _0241_ ;
wire _0242_ ;
wire _0243_ ;
wire _0244_ ;
wire _0245_ ;
wire _0246_ ;
wire _0247_ ;
wire _0248_ ;
wire _0249_ ;
wire _0250_ ;
wire _0251_ ;
wire _0252_ ;
wire _0253_ ;
wire _0254_ ;
wire _0255_ ;
wire _0256_ ;
wire _0257_ ;
wire _0258_ ;
wire _0259_ ;
wire _0260_ ;
wire _0261_ ;
wire _0262_ ;
wire _0263_ ;
wire _0264_ ;
wire _0265_ ;
wire _0266_ ;
wire _0267_ ;
wire _0268_ ;
wire _0269_ ;
wire _0270_ ;
wire _0271_ ;
wire _0272_ ;
wire _0273_ ;
wire _0274_ ;
wire _0275_ ;
wire _0276_ ;
wire _0277_ ;
wire _0278_ ;
wire _0279_ ;
wire _0280_ ;
wire _0281_ ;
wire _0282_ ;
wire _0283_ ;
wire _0284_ ;
wire _0285_ ;
wire _0286_ ;
wire _0287_ ;
wire _0288_ ;
wire _0289_ ;
wire _0290_ ;
wire _0291_ ;
wire _0292_ ;
wire _0293_ ;
wire _0294_ ;
wire _0295_ ;
wire _0296_ ;
wire _0297_ ;
wire _0298_ ;
wire _0299_ ;
wire _0300_ ;
wire _0301_ ;
wire _0302_ ;
wire _0303_ ;
wire _0304_ ;
wire _0305_ ;
wire _0306_ ;
wire _0307_ ;
wire _0308_ ;
wire _0309_ ;
wire _0310_ ;
wire _0311_ ;
wire _0312_ ;
wire _0313_ ;
wire _0314_ ;
wire _0315_ ;
wire _0316_ ;
wire _0317_ ;
wire _0318_ ;
wire _0319_ ;
wire _0320_ ;
wire _0321_ ;
wire _0322_ ;
wire _0323_ ;
wire _0324_ ;
wire _0325_ ;
wire _0326_ ;
wire _0327_ ;
wire _0328_ ;
wire _0329_ ;
wire _0330_ ;
wire _0331_ ;
wire _0332_ ;
wire _0333_ ;
wire _0334_ ;
wire _0335_ ;
wire _0336_ ;
wire _0337_ ;
wire _0338_ ;
wire _0339_ ;
wire _0340_ ;
wire _0341_ ;
wire _0342_ ;
wire _0343_ ;
wire _0344_ ;
wire _0345_ ;
wire _0346_ ;
wire _0347_ ;
wire _0348_ ;
wire _0349_ ;
wire _0350_ ;
wire _0351_ ;
wire _0352_ ;
wire _0353_ ;
wire _0354_ ;
wire _0355_ ;
wire _0356_ ;
wire _0357_ ;
wire _0358_ ;
wire _0359_ ;
wire _0360_ ;
wire _0361_ ;
wire _0362_ ;
wire _0363_ ;
wire _0364_ ;
wire _0365_ ;
wire _0366_ ;
wire _0367_ ;
wire _0368_ ;
wire _0369_ ;
wire _0370_ ;
wire _0371_ ;
wire _0372_ ;
wire _0373_ ;
wire _0374_ ;
wire _0375_ ;
wire _0376_ ;
wire _0377_ ;
wire _0378_ ;
wire _0379_ ;
wire _0380_ ;
wire _0381_ ;
wire _0382_ ;
wire _0383_ ;
wire _0384_ ;
wire _0385_ ;
wire _0386_ ;
wire _0387_ ;
wire _0388_ ;
wire _0389_ ;
wire _0390_ ;
wire _0391_ ;
wire _0392_ ;
wire _0393_ ;
wire _0394_ ;
wire _0395_ ;
wire _0396_ ;
wire _0397_ ;
wire _0398_ ;
wire _0399_ ;
wire _0400_ ;
wire _0401_ ;
wire _0402_ ;
wire _0403_ ;
wire _0404_ ;
wire _0405_ ;
wire _0406_ ;
wire _0407_ ;
wire _0408_ ;
wire _0409_ ;
wire _0410_ ;
wire _0411_ ;
wire _0412_ ;
wire _0413_ ;
wire _0414_ ;
wire _0415_ ;
wire _0416_ ;
wire _0417_ ;
wire _0418_ ;
wire _0419_ ;
wire _0420_ ;
wire _0421_ ;
wire _0422_ ;
wire _0423_ ;
wire _0424_ ;
wire _0425_ ;
wire _0426_ ;
wire _0427_ ;
wire _0428_ ;
wire _0429_ ;
wire _0430_ ;
wire _0431_ ;
wire _0432_ ;
wire _0433_ ;
wire _0434_ ;
wire _0435_ ;
wire _0436_ ;
wire _0437_ ;
wire _0438_ ;
wire _0439_ ;
wire _0440_ ;
wire _0441_ ;
wire _0442_ ;
wire _0443_ ;
wire _0444_ ;
wire _0445_ ;
wire _0446_ ;
wire _0447_ ;
wire _0448_ ;
wire _0449_ ;
wire _0450_ ;
wire _0451_ ;
wire _0452_ ;
wire _0453_ ;
wire _0454_ ;
wire _0455_ ;
wire _0456_ ;
wire _0457_ ;
wire _0458_ ;
wire _0459_ ;
wire _0460_ ;
wire _0461_ ;
wire _0462_ ;
wire _0463_ ;
wire _0464_ ;
wire _0465_ ;
wire _0466_ ;
wire _0467_ ;
wire _0468_ ;
wire _0469_ ;
wire _0470_ ;
wire _0471_ ;
wire _0472_ ;
wire _0473_ ;
wire _0474_ ;
wire _0475_ ;
wire _0476_ ;
wire _0477_ ;
wire _0478_ ;
wire _0479_ ;
wire _0480_ ;
wire _0481_ ;
wire _0482_ ;
wire _0483_ ;
wire _0484_ ;
wire _0485_ ;
wire _0486_ ;
wire _0487_ ;
wire _0488_ ;
wire _0489_ ;
wire _0490_ ;
wire _0491_ ;
wire _0492_ ;
wire _0493_ ;
wire _0494_ ;
wire _0495_ ;
wire _0496_ ;
wire _0497_ ;
wire _0498_ ;
wire _0499_ ;
wire _0500_ ;
wire _0501_ ;
wire _0502_ ;
wire _0503_ ;
wire _0504_ ;
wire _0505_ ;
wire _0506_ ;
wire _0507_ ;
wire _0508_ ;
wire _0509_ ;
wire _0510_ ;
wire _0511_ ;
wire _0512_ ;
wire _0513_ ;
wire _0514_ ;
wire _0515_ ;
wire _0516_ ;
wire _0517_ ;
wire _0518_ ;
wire _0519_ ;
wire _0520_ ;
wire _0521_ ;
wire _0522_ ;
wire _0523_ ;
wire _0524_ ;
wire _0525_ ;
wire _0526_ ;
wire _0527_ ;
wire _0528_ ;
wire _0529_ ;
wire _0530_ ;
wire _0531_ ;
wire _0532_ ;
wire _0533_ ;
wire _0534_ ;
wire _0535_ ;
wire _0536_ ;
wire _0537_ ;
wire _0538_ ;
wire _0539_ ;
wire _0540_ ;
wire _0541_ ;
wire _0542_ ;
wire _0543_ ;
wire _0544_ ;
wire _0545_ ;
wire _0546_ ;
wire _0547_ ;
wire _0548_ ;
wire _0549_ ;
wire _0550_ ;
wire _0551_ ;
wire _0552_ ;
wire _0553_ ;
wire _0554_ ;
wire _0555_ ;
wire _0556_ ;
wire _0557_ ;
wire _0558_ ;
wire _0559_ ;
wire _0560_ ;
wire _0561_ ;
wire _0562_ ;
wire _0563_ ;
wire _0564_ ;
wire _0565_ ;
wire _0566_ ;
wire _0567_ ;
wire _0568_ ;
wire _0569_ ;
wire _0570_ ;
wire _0571_ ;
wire _0572_ ;
wire _0573_ ;
wire _0574_ ;
wire _0575_ ;
wire _0576_ ;
wire _0577_ ;
wire _0578_ ;
wire _0579_ ;
wire _0580_ ;
wire _0581_ ;
wire _0582_ ;
wire _0583_ ;
wire _0584_ ;
wire _0585_ ;
wire _0586_ ;
wire _0587_ ;
wire _0588_ ;
wire _0589_ ;
wire _0590_ ;
wire _0591_ ;
wire _0592_ ;
wire _0593_ ;
wire _0594_ ;
wire _0595_ ;
wire _0596_ ;
wire _0597_ ;
wire _0598_ ;
wire _0599_ ;
wire _0600_ ;
wire _0601_ ;
wire _0602_ ;
wire _0603_ ;
wire _0604_ ;
wire _0605_ ;
wire _0606_ ;
wire _0607_ ;
wire _0608_ ;
wire _0609_ ;
wire _0610_ ;
wire _0611_ ;
wire _0612_ ;
wire _0613_ ;
wire _0614_ ;
wire _0615_ ;
wire _0616_ ;
wire _0617_ ;
wire _0618_ ;
wire _0619_ ;
wire _0620_ ;
wire _0621_ ;
wire _0622_ ;
wire _0623_ ;
wire _0624_ ;
wire _0625_ ;
wire _0626_ ;
wire _0627_ ;
wire _0628_ ;
wire _0629_ ;
wire _0630_ ;
wire _0631_ ;
wire _0632_ ;
wire _0633_ ;
wire _0634_ ;
wire _0635_ ;
wire _0636_ ;
wire _0637_ ;
wire _0638_ ;
wire _0639_ ;
wire _0640_ ;
wire _0641_ ;
wire _0642_ ;
wire _0643_ ;
wire _0644_ ;
wire _0645_ ;
wire _0646_ ;
wire _0647_ ;
wire _0648_ ;
wire _0649_ ;
wire _0650_ ;
wire _0651_ ;
wire _0652_ ;
wire _0653_ ;
wire _0654_ ;
wire _0655_ ;
wire _0656_ ;
wire _0657_ ;
wire _0658_ ;
wire _0659_ ;
wire _0660_ ;
wire _0661_ ;
wire _0662_ ;
wire _0663_ ;
wire _0664_ ;
wire _0665_ ;
wire _0666_ ;
wire _0667_ ;
wire _0668_ ;
wire _0669_ ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire \b[0] ;
wire \b[1] ;
wire \b[2] ;
wire \b[3] ;
wire \b[4] ;
wire \b[5] ;
wire \b[6] ;
wire \b[7] ;
wire \b[8] ;
wire \b[9] ;
wire \b[10] ;
wire \b[11] ;
wire \b[12] ;
wire \b[13] ;
wire \b[14] ;
wire \b[15] ;
wire \b[16] ;
wire \b[17] ;
wire \b[18] ;
wire \b[19] ;
wire \b[20] ;
wire \b[21] ;
wire \b[22] ;
wire \b[23] ;
wire \b[24] ;
wire \b[25] ;
wire \b[26] ;
wire \b[27] ;
wire \b[28] ;
wire \b[29] ;
wire \b[30] ;
wire \b[31] ;
wire \a[0] ;
wire \a[1] ;
wire \a[2] ;
wire \a[3] ;
wire \a[4] ;
wire \a[5] ;
wire \a[6] ;
wire \a[7] ;
wire \a[8] ;
wire \a[9] ;
wire \a[10] ;
wire \a[11] ;
wire \a[12] ;
wire \a[13] ;
wire \a[14] ;
wire \a[15] ;
wire \a[16] ;
wire \a[17] ;
wire \a[18] ;
wire \a[19] ;
wire \a[20] ;
wire \a[21] ;
wire \a[22] ;
wire \a[23] ;
wire \a[24] ;
wire \a[25] ;
wire \a[26] ;
wire \a[27] ;
wire \a[28] ;
wire \a[29] ;
wire \a[30] ;
wire \a[31] ;
wire \ctrl[0] ;
wire \ctrl[1] ;
wire \ctrl[2] ;
wire \ctrl[3] ;
wire \result[0] ;
wire \result[1] ;
wire \result[2] ;
wire \result[3] ;
wire \result[4] ;
wire \result[5] ;
wire \result[6] ;
wire \result[7] ;
wire \result[8] ;
wire \result[9] ;
wire \result[10] ;
wire \result[11] ;
wire \result[12] ;
wire \result[13] ;
wire \result[14] ;
wire \result[15] ;
wire \result[16] ;
wire \result[17] ;
wire \result[18] ;
wire \result[19] ;
wire \result[20] ;
wire \result[21] ;
wire \result[22] ;
wire \result[23] ;
wire \result[24] ;
wire \result[25] ;
wire \result[26] ;
wire \result[27] ;
wire \result[28] ;
wire \result[29] ;
wire \result[30] ;
wire \result[31] ;

assign \b[0] = b[0] ;
assign \b[1] = b[1] ;
assign \b[2] = b[2] ;
assign \b[3] = b[3] ;
assign \b[4] = b[4] ;
assign \a[0] = a[0] ;
assign \a[1] = a[1] ;
assign \a[2] = a[2] ;
assign \a[3] = a[3] ;
assign \a[4] = a[4] ;
assign \a[5] = a[5] ;
assign \a[6] = a[6] ;
assign \a[7] = a[7] ;
assign \a[8] = a[8] ;
assign \a[9] = a[9] ;
assign \a[10] = a[10] ;
assign \a[11] = a[11] ;
assign \a[12] = a[12] ;
assign \a[13] = a[13] ;
assign \a[14] = a[14] ;
assign \a[15] = a[15] ;
assign \a[16] = a[16] ;
assign \a[17] = a[17] ;
assign \a[18] = a[18] ;
assign \a[19] = a[19] ;
assign \a[20] = a[20] ;
assign \a[21] = a[21] ;
assign \a[22] = a[22] ;
assign \a[23] = a[23] ;
assign \a[24] = a[24] ;
assign \a[25] = a[25] ;
assign \a[26] = a[26] ;
assign \a[27] = a[27] ;
assign \a[28] = a[28] ;
assign \a[29] = a[29] ;
assign \a[30] = a[30] ;
assign \a[31] = a[31] ;
assign \ctrl[0] = ctrl[0] ;
assign \ctrl[1] = ctrl[1] ;
assign \ctrl[2] = ctrl[2] ;
assign \ctrl[3] = ctrl[3] ;
assign result[0] = \result[0] ;
assign result[1] = \result[1] ;
assign result[2] = \result[2] ;
assign result[3] = \result[3] ;
assign result[4] = \result[4] ;
assign result[5] = \result[5] ;
assign result[6] = \result[6] ;
assign result[7] = \result[7] ;
assign result[8] = \result[8] ;
assign result[9] = \result[9] ;
assign result[10] = \result[10] ;
assign result[11] = \result[11] ;
assign result[12] = \result[12] ;
assign result[13] = \result[13] ;
assign result[14] = \result[14] ;
assign result[15] = \result[15] ;
assign result[16] = \result[16] ;
assign result[17] = \result[17] ;
assign result[18] = \result[18] ;
assign result[19] = \result[19] ;
assign result[20] = \result[20] ;
assign result[21] = \result[21] ;
assign result[22] = \result[22] ;
assign result[23] = \result[23] ;
assign result[24] = \result[24] ;
assign result[25] = \result[25] ;
assign result[26] = \result[26] ;
assign result[27] = \result[27] ;
assign result[28] = \result[28] ;
assign result[29] = \result[29] ;
assign result[30] = \result[30] ;
assign result[31] = \result[31] ;

NOR2_X1 _0670_ ( .A1(fanout_net_1 ), .A2(_0016_ ), .ZN(_0612_ ) );
INV_X1 _0671_ ( .A(_0612_ ), .ZN(_0613_ ) );
INV_X32 _0672_ ( .A(fanout_net_2 ), .ZN(_0614_ ) );
BUF_X32 _0673_ ( .A(_0614_ ), .Z(_0615_ ) );
BUF_X4 _0674_ ( .A(_0615_ ), .Z(_0616_ ) );
INV_X32 _0675_ ( .A(fanout_net_1 ), .ZN(_0617_ ) );
BUF_X32 _0676_ ( .A(_0617_ ), .Z(_0618_ ) );
BUF_X32 _0677_ ( .A(_0618_ ), .Z(_0619_ ) );
OAI211_X2 _0678_ ( .A(_0613_ ), .B(_0616_ ), .C1(_0619_ ), .C2(_0017_ ), .ZN(_0620_ ) );
NOR2_X1 _0679_ ( .A1(fanout_net_1 ), .A2(_0018_ ), .ZN(_0621_ ) );
INV_X1 _0680_ ( .A(_0621_ ), .ZN(_0622_ ) );
OAI211_X2 _0681_ ( .A(_0622_ ), .B(fanout_net_2 ), .C1(_0619_ ), .C2(_0019_ ), .ZN(_0623_ ) );
INV_X1 _0682_ ( .A(fanout_net_4 ), .ZN(_0624_ ) );
BUF_X2 _0683_ ( .A(_0624_ ), .Z(_0625_ ) );
NAND3_X1 _0684_ ( .A1(_0620_ ), .A2(_0623_ ), .A3(_0625_ ), .ZN(_0626_ ) );
NOR2_X1 _0685_ ( .A1(fanout_net_1 ), .A2(_0023_ ), .ZN(_0627_ ) );
INV_X1 _0686_ ( .A(_0024_ ), .ZN(_0628_ ) );
AOI21_X1 _0687_ ( .A(_0627_ ), .B1(fanout_net_1 ), .B2(_0628_ ), .ZN(_0629_ ) );
BUF_X32 _0688_ ( .A(_0618_ ), .Z(_0630_ ) );
NOR2_X4 _0689_ ( .A1(_0630_ ), .A2(_0021_ ), .ZN(_0631_ ) );
NOR2_X1 _0690_ ( .A1(fanout_net_1 ), .A2(_0020_ ), .ZN(_0632_ ) );
NOR2_X1 _0691_ ( .A1(_0631_ ), .A2(_0632_ ), .ZN(_0633_ ) );
MUX2_X2 _0692_ ( .A(_0629_ ), .B(_0633_ ), .S(_0616_ ), .Z(_0634_ ) );
BUF_X4 _0693_ ( .A(_0624_ ), .Z(_0635_ ) );
BUF_X4 _0694_ ( .A(_0635_ ), .Z(_0636_ ) );
OAI21_X2 _0695_ ( .A(_0626_ ), .B1(_0634_ ), .B2(_0636_ ), .ZN(_0637_ ) );
INV_X1 _0696_ ( .A(fanout_net_6 ), .ZN(_0041_ ) );
BUF_X4 _0697_ ( .A(_0041_ ), .Z(_0042_ ) );
NOR2_X1 _0698_ ( .A1(_0637_ ), .A2(_0042_ ), .ZN(_0043_ ) );
NOR2_X1 _0699_ ( .A1(_0617_ ), .A2(_0010_ ), .ZN(_0044_ ) );
NOR2_X1 _0700_ ( .A1(fanout_net_1 ), .A2(_0009_ ), .ZN(_0045_ ) );
NOR3_X1 _0701_ ( .A1(_0044_ ), .A2(_0615_ ), .A3(_0045_ ), .ZN(_0046_ ) );
NOR2_X4 _0702_ ( .A1(_0618_ ), .A2(_0008_ ), .ZN(_0047_ ) );
NOR2_X1 _0703_ ( .A1(fanout_net_1 ), .A2(_0007_ ), .ZN(_0048_ ) );
NOR3_X1 _0704_ ( .A1(_0047_ ), .A2(fanout_net_2 ), .A3(_0048_ ), .ZN(_0049_ ) );
NOR2_X1 _0705_ ( .A1(_0046_ ), .A2(_0049_ ), .ZN(_0050_ ) );
NAND2_X1 _0706_ ( .A1(_0050_ ), .A2(_0625_ ), .ZN(_0051_ ) );
NOR2_X4 _0707_ ( .A1(_0630_ ), .A2(_0015_ ), .ZN(_0052_ ) );
NOR2_X1 _0708_ ( .A1(fanout_net_1 ), .A2(_0014_ ), .ZN(_0053_ ) );
NOR3_X1 _0709_ ( .A1(_0052_ ), .A2(_0615_ ), .A3(_0053_ ), .ZN(_0054_ ) );
NOR2_X2 _0710_ ( .A1(_0618_ ), .A2(_0013_ ), .ZN(_0055_ ) );
NOR2_X1 _0711_ ( .A1(fanout_net_1 ), .A2(_0012_ ), .ZN(_0056_ ) );
NOR3_X1 _0712_ ( .A1(_0055_ ), .A2(fanout_net_2 ), .A3(_0056_ ), .ZN(_0057_ ) );
NOR2_X1 _0713_ ( .A1(_0054_ ), .A2(_0057_ ), .ZN(_0058_ ) );
NAND2_X1 _0714_ ( .A1(_0058_ ), .A2(fanout_net_4 ), .ZN(_0059_ ) );
BUF_X2 _0715_ ( .A(_0041_ ), .Z(_0060_ ) );
AND3_X1 _0716_ ( .A1(_0051_ ), .A2(_0059_ ), .A3(_0060_ ), .ZN(_0061_ ) );
INV_X1 _0717_ ( .A(fanout_net_7 ), .ZN(_0062_ ) );
BUF_X4 _0718_ ( .A(_0062_ ), .Z(_0063_ ) );
OR3_X2 _0719_ ( .A1(_0043_ ), .A2(_0061_ ), .A3(_0063_ ), .ZN(_0064_ ) );
INV_X1 _0720_ ( .A(_0037_ ), .ZN(_0065_ ) );
NOR2_X1 _0721_ ( .A1(_0065_ ), .A2(_0038_ ), .ZN(_0066_ ) );
INV_X1 _0722_ ( .A(_0039_ ), .ZN(_0067_ ) );
NOR2_X1 _0723_ ( .A1(_0067_ ), .A2(_0040_ ), .ZN(_0068_ ) );
AND2_X1 _0724_ ( .A1(_0066_ ), .A2(_0068_ ), .ZN(_0069_ ) );
BUF_X4 _0725_ ( .A(_0069_ ), .Z(_0070_ ) );
BUF_X4 _0726_ ( .A(_0063_ ), .Z(_0071_ ) );
NOR2_X1 _0727_ ( .A1(_0619_ ), .A2(_0029_ ), .ZN(_0072_ ) );
NOR2_X1 _0728_ ( .A1(fanout_net_1 ), .A2(_0028_ ), .ZN(_0073_ ) );
OAI21_X1 _0729_ ( .A(fanout_net_2 ), .B1(_0072_ ), .B2(_0073_ ), .ZN(_0074_ ) );
NAND2_X1 _0730_ ( .A1(_0619_ ), .A2(_0026_ ), .ZN(_0075_ ) );
BUF_X16 _0731_ ( .A(_0615_ ), .Z(_0076_ ) );
BUF_X32 _0732_ ( .A(_0630_ ), .Z(_0077_ ) );
INV_X1 _0733_ ( .A(_0027_ ), .ZN(_0078_ ) );
OAI211_X2 _0734_ ( .A(_0075_ ), .B(_0076_ ), .C1(_0077_ ), .C2(_0078_ ), .ZN(_0079_ ) );
AND3_X1 _0735_ ( .A1(_0074_ ), .A2(_0079_ ), .A3(fanout_net_4 ), .ZN(_0080_ ) );
MUX2_X1 _0736_ ( .A(_0000_ ), .B(_0011_ ), .S(fanout_net_1 ), .Z(_0081_ ) );
INV_X1 _0737_ ( .A(_0022_ ), .ZN(_0082_ ) );
NOR2_X1 _0738_ ( .A1(_0082_ ), .A2(fanout_net_1 ), .ZN(_0083_ ) );
INV_X1 _0739_ ( .A(_0083_ ), .ZN(_0084_ ) );
NAND2_X1 _0740_ ( .A1(fanout_net_1 ), .A2(_0025_ ), .ZN(_0085_ ) );
NAND2_X1 _0741_ ( .A1(_0084_ ), .A2(_0085_ ), .ZN(_0086_ ) );
MUX2_X1 _0742_ ( .A(_0081_ ), .B(_0086_ ), .S(fanout_net_2 ), .Z(_0087_ ) );
BUF_X4 _0743_ ( .A(_0635_ ), .Z(_0088_ ) );
AOI211_X2 _0744_ ( .A(fanout_net_6 ), .B(_0080_ ), .C1(_0087_ ), .C2(_0088_ ), .ZN(_0089_ ) );
NOR2_X1 _0745_ ( .A1(fanout_net_1 ), .A2(_0005_ ), .ZN(_0090_ ) );
INV_X1 _0746_ ( .A(_0090_ ), .ZN(_0091_ ) );
OAI211_X2 _0747_ ( .A(_0091_ ), .B(fanout_net_2 ), .C1(_0077_ ), .C2(_0006_ ), .ZN(_0092_ ) );
NOR2_X1 _0748_ ( .A1(fanout_net_1 ), .A2(_0003_ ), .ZN(_0093_ ) );
INV_X1 _0749_ ( .A(_0093_ ), .ZN(_0094_ ) );
OAI211_X2 _0750_ ( .A(_0094_ ), .B(_0616_ ), .C1(_0077_ ), .C2(_0004_ ), .ZN(_0095_ ) );
AND3_X1 _0751_ ( .A1(_0092_ ), .A2(_0095_ ), .A3(fanout_net_4 ), .ZN(_0096_ ) );
BUF_X4 _0752_ ( .A(_0076_ ), .Z(_0097_ ) );
NOR2_X4 _0753_ ( .A1(_0619_ ), .A2(_0031_ ), .ZN(_0098_ ) );
NOR2_X1 _0754_ ( .A1(fanout_net_1 ), .A2(_0030_ ), .ZN(_0099_ ) );
OAI21_X1 _0755_ ( .A(_0097_ ), .B1(_0098_ ), .B2(_0099_ ), .ZN(_0100_ ) );
NOR2_X4 _0756_ ( .A1(_0630_ ), .A2(_0002_ ), .ZN(_0101_ ) );
NOR2_X1 _0757_ ( .A1(fanout_net_1 ), .A2(_0001_ ), .ZN(_0102_ ) );
OAI21_X1 _0758_ ( .A(fanout_net_2 ), .B1(_0101_ ), .B2(_0102_ ), .ZN(_0103_ ) );
AOI21_X1 _0759_ ( .A(fanout_net_4 ), .B1(_0100_ ), .B2(_0103_ ), .ZN(_0104_ ) );
NOR2_X1 _0760_ ( .A1(_0096_ ), .A2(_0104_ ), .ZN(_0105_ ) );
BUF_X2 _0761_ ( .A(_0060_ ), .Z(_0106_ ) );
NOR2_X1 _0762_ ( .A1(_0105_ ), .A2(_0106_ ), .ZN(_0107_ ) );
OAI21_X1 _0763_ ( .A(_0071_ ), .B1(_0089_ ), .B2(_0107_ ), .ZN(_0108_ ) );
NAND3_X1 _0764_ ( .A1(_0064_ ), .A2(_0070_ ), .A3(_0108_ ), .ZN(_0109_ ) );
OR3_X1 _0765_ ( .A1(_0065_ ), .A2(_0038_ ), .A3(_0039_ ), .ZN(_0110_ ) );
NOR2_X4 _0766_ ( .A1(_0110_ ), .A2(_0040_ ), .ZN(_0111_ ) );
BUF_X4 _0767_ ( .A(_0111_ ), .Z(_0112_ ) );
BUF_X4 _0768_ ( .A(_0106_ ), .Z(_0113_ ) );
INV_X1 _0769_ ( .A(_0000_ ), .ZN(_0114_ ) );
NOR2_X1 _0770_ ( .A1(_0114_ ), .A2(fanout_net_1 ), .ZN(_0115_ ) );
AND3_X1 _0771_ ( .A1(_0115_ ), .A2(_0635_ ), .A3(_0097_ ), .ZN(_0116_ ) );
NAND4_X1 _0772_ ( .A1(_0112_ ), .A2(_0113_ ), .A3(_0071_ ), .A4(_0116_ ), .ZN(_0117_ ) );
NAND2_X1 _0773_ ( .A1(_0109_ ), .A2(_0117_ ), .ZN(_0638_ ) );
NOR2_X1 _0774_ ( .A1(_0630_ ), .A2(_0018_ ), .ZN(_0118_ ) );
NOR2_X1 _0775_ ( .A1(fanout_net_1 ), .A2(_0017_ ), .ZN(_0119_ ) );
OAI21_X1 _0776_ ( .A(_0076_ ), .B1(_0118_ ), .B2(_0119_ ), .ZN(_0120_ ) );
NOR2_X4 _0777_ ( .A1(_0630_ ), .A2(_0020_ ), .ZN(_0121_ ) );
NOR2_X1 _0778_ ( .A1(fanout_net_1 ), .A2(_0019_ ), .ZN(_0122_ ) );
OAI21_X1 _0779_ ( .A(fanout_net_2 ), .B1(_0121_ ), .B2(_0122_ ), .ZN(_0123_ ) );
NAND2_X1 _0780_ ( .A1(_0120_ ), .A2(_0123_ ), .ZN(_0124_ ) );
OR2_X4 _0781_ ( .A1(_0630_ ), .A2(_0023_ ), .ZN(_0125_ ) );
NOR2_X1 _0782_ ( .A1(fanout_net_1 ), .A2(_0021_ ), .ZN(_0126_ ) );
INV_X1 _0783_ ( .A(_0126_ ), .ZN(_0127_ ) );
NAND2_X4 _0784_ ( .A1(_0125_ ), .A2(_0127_ ), .ZN(_0128_ ) );
NAND2_X1 _0785_ ( .A1(_0128_ ), .A2(_0076_ ), .ZN(_0129_ ) );
BUF_X4 _0786_ ( .A(_0615_ ), .Z(_0130_ ) );
NOR2_X1 _0787_ ( .A1(_0628_ ), .A2(fanout_net_1 ), .ZN(_0131_ ) );
OAI21_X2 _0788_ ( .A(_0129_ ), .B1(_0130_ ), .B2(_0131_ ), .ZN(_0132_ ) );
MUX2_X2 _0789_ ( .A(_0124_ ), .B(_0132_ ), .S(fanout_net_4 ), .Z(_0133_ ) );
NOR2_X1 _0790_ ( .A1(_0133_ ), .A2(_0042_ ), .ZN(_0134_ ) );
NOR2_X4 _0791_ ( .A1(_0630_ ), .A2(_0016_ ), .ZN(_0135_ ) );
NOR2_X1 _0792_ ( .A1(fanout_net_1 ), .A2(_0015_ ), .ZN(_0136_ ) );
NOR3_X1 _0793_ ( .A1(_0135_ ), .A2(_0616_ ), .A3(_0136_ ), .ZN(_0137_ ) );
NOR2_X1 _0794_ ( .A1(_0617_ ), .A2(_0014_ ), .ZN(_0138_ ) );
NOR2_X1 _0795_ ( .A1(fanout_net_1 ), .A2(_0013_ ), .ZN(_0139_ ) );
NOR3_X1 _0796_ ( .A1(_0138_ ), .A2(fanout_net_2 ), .A3(_0139_ ), .ZN(_0140_ ) );
NOR2_X1 _0797_ ( .A1(_0137_ ), .A2(_0140_ ), .ZN(_0141_ ) );
NAND2_X1 _0798_ ( .A1(_0141_ ), .A2(fanout_net_4 ), .ZN(_0142_ ) );
NOR2_X4 _0799_ ( .A1(_0619_ ), .A2(_0009_ ), .ZN(_0143_ ) );
NOR2_X4 _0800_ ( .A1(fanout_net_1 ), .A2(_0008_ ), .ZN(_0144_ ) );
OAI21_X1 _0801_ ( .A(_0076_ ), .B1(_0143_ ), .B2(_0144_ ), .ZN(_0145_ ) );
NOR2_X1 _0802_ ( .A1(_0617_ ), .A2(_0012_ ), .ZN(_0146_ ) );
NOR2_X1 _0803_ ( .A1(fanout_net_1 ), .A2(_0010_ ), .ZN(_0147_ ) );
OAI21_X1 _0804_ ( .A(fanout_net_2 ), .B1(_0146_ ), .B2(_0147_ ), .ZN(_0148_ ) );
NAND2_X1 _0805_ ( .A1(_0145_ ), .A2(_0148_ ), .ZN(_0149_ ) );
NAND2_X1 _0806_ ( .A1(_0149_ ), .A2(_0625_ ), .ZN(_0150_ ) );
AND3_X1 _0807_ ( .A1(_0142_ ), .A2(_0060_ ), .A3(_0150_ ), .ZN(_0151_ ) );
OR3_X4 _0808_ ( .A1(_0134_ ), .A2(_0063_ ), .A3(_0151_ ), .ZN(_0152_ ) );
BUF_X2 _0809_ ( .A(_0042_ ), .Z(_0153_ ) );
NOR2_X1 _0810_ ( .A1(_0011_ ), .A2(fanout_net_1 ), .ZN(_0154_ ) );
AOI21_X1 _0811_ ( .A(_0154_ ), .B1(fanout_net_1 ), .B2(_0082_ ), .ZN(_0155_ ) );
NOR2_X1 _0812_ ( .A1(_0155_ ), .A2(fanout_net_2 ), .ZN(_0156_ ) );
NOR2_X4 _0813_ ( .A1(_0077_ ), .A2(_0026_ ), .ZN(_0157_ ) );
NOR2_X1 _0814_ ( .A1(fanout_net_1 ), .A2(_0025_ ), .ZN(_0158_ ) );
OR2_X1 _0815_ ( .A1(_0157_ ), .A2(_0158_ ), .ZN(_0159_ ) );
AOI211_X2 _0816_ ( .A(fanout_net_4 ), .B(_0156_ ), .C1(fanout_net_2 ), .C2(_0159_ ), .ZN(_0160_ ) );
BUF_X4 _0817_ ( .A(_0636_ ), .Z(_0161_ ) );
NOR2_X1 _0818_ ( .A1(_0032_ ), .A2(_0029_ ), .ZN(_0162_ ) );
INV_X1 _0819_ ( .A(_0162_ ), .ZN(_0163_ ) );
BUF_X32 _0820_ ( .A(_0077_ ), .Z(_0164_ ) );
OAI211_X2 _0821_ ( .A(_0163_ ), .B(fanout_net_2 ), .C1(_0164_ ), .C2(_0030_ ), .ZN(_0165_ ) );
NOR2_X1 _0822_ ( .A1(_0032_ ), .A2(_0027_ ), .ZN(_0166_ ) );
INV_X1 _0823_ ( .A(_0166_ ), .ZN(_0167_ ) );
BUF_X4 _0824_ ( .A(_0130_ ), .Z(_0168_ ) );
OAI211_X2 _0825_ ( .A(_0167_ ), .B(_0168_ ), .C1(_0164_ ), .C2(_0028_ ), .ZN(_0169_ ) );
AOI21_X1 _0826_ ( .A(_0161_ ), .B1(_0165_ ), .B2(_0169_ ), .ZN(_0170_ ) );
OAI21_X1 _0827_ ( .A(_0153_ ), .B1(_0160_ ), .B2(_0170_ ), .ZN(_0171_ ) );
NOR2_X1 _0828_ ( .A1(_0032_ ), .A2(_0006_ ), .ZN(_0172_ ) );
INV_X1 _0829_ ( .A(_0172_ ), .ZN(_0173_ ) );
OAI211_X2 _0830_ ( .A(_0173_ ), .B(fanout_net_2 ), .C1(_0619_ ), .C2(_0007_ ), .ZN(_0174_ ) );
NOR2_X1 _0831_ ( .A1(_0032_ ), .A2(_0004_ ), .ZN(_0175_ ) );
INV_X1 _0832_ ( .A(_0175_ ), .ZN(_0176_ ) );
OAI211_X2 _0833_ ( .A(_0176_ ), .B(_0615_ ), .C1(_0619_ ), .C2(_0005_ ), .ZN(_0177_ ) );
AOI21_X1 _0834_ ( .A(_0636_ ), .B1(_0174_ ), .B2(_0177_ ), .ZN(_0178_ ) );
NOR2_X1 _0835_ ( .A1(_0618_ ), .A2(_0001_ ), .ZN(_0179_ ) );
NOR2_X1 _0836_ ( .A1(_0032_ ), .A2(_0031_ ), .ZN(_0180_ ) );
OAI21_X1 _0837_ ( .A(_0097_ ), .B1(_0179_ ), .B2(_0180_ ), .ZN(_0181_ ) );
NOR2_X1 _0838_ ( .A1(_0618_ ), .A2(_0003_ ), .ZN(_0182_ ) );
NOR2_X1 _0839_ ( .A1(_0032_ ), .A2(_0002_ ), .ZN(_0183_ ) );
OAI21_X1 _0840_ ( .A(fanout_net_2 ), .B1(_0182_ ), .B2(_0183_ ), .ZN(_0184_ ) );
AND3_X1 _0841_ ( .A1(_0181_ ), .A2(_0184_ ), .A3(_0636_ ), .ZN(_0185_ ) );
OAI21_X1 _0842_ ( .A(fanout_net_6 ), .B1(_0178_ ), .B2(_0185_ ), .ZN(_0186_ ) );
NAND3_X1 _0843_ ( .A1(_0171_ ), .A2(_0071_ ), .A3(_0186_ ), .ZN(_0187_ ) );
NAND3_X1 _0844_ ( .A1(_0152_ ), .A2(_0070_ ), .A3(_0187_ ), .ZN(_0188_ ) );
AOI21_X1 _0845_ ( .A(_0154_ ), .B1(_0114_ ), .B2(_0032_ ), .ZN(_0189_ ) );
AND3_X1 _0846_ ( .A1(_0189_ ), .A2(_0088_ ), .A3(_0168_ ), .ZN(_0190_ ) );
NAND4_X1 _0847_ ( .A1(_0190_ ), .A2(_0113_ ), .A3(_0071_ ), .A4(_0112_ ), .ZN(_0191_ ) );
NAND2_X1 _0848_ ( .A1(_0188_ ), .A2(_0191_ ), .ZN(_0649_ ) );
AND2_X2 _0849_ ( .A1(_0111_ ), .A2(_0063_ ), .ZN(_0192_ ) );
AND2_X1 _0850_ ( .A1(_0011_ ), .A2(_0032_ ), .ZN(_0193_ ) );
OAI21_X1 _0851_ ( .A(_0130_ ), .B1(_0083_ ), .B2(_0193_ ), .ZN(_0194_ ) );
NAND3_X1 _0852_ ( .A1(_0164_ ), .A2(fanout_net_2 ), .A3(_0000_ ), .ZN(_0195_ ) );
AOI21_X1 _0853_ ( .A(fanout_net_4 ), .B1(_0194_ ), .B2(_0195_ ), .ZN(_0196_ ) );
NAND3_X1 _0854_ ( .A1(_0192_ ), .A2(_0113_ ), .A3(_0196_ ), .ZN(_0197_ ) );
BUF_X2 _0855_ ( .A(_0042_ ), .Z(_0198_ ) );
NOR2_X4 _0856_ ( .A1(_0630_ ), .A2(_0004_ ), .ZN(_0199_ ) );
BUF_X4 _0857_ ( .A(_0130_ ), .Z(_0200_ ) );
NOR3_X1 _0858_ ( .A1(_0199_ ), .A2(_0200_ ), .A3(_0093_ ), .ZN(_0201_ ) );
NOR3_X1 _0859_ ( .A1(_0101_ ), .A2(fanout_net_2 ), .A3(_0102_ ), .ZN(_0202_ ) );
NOR2_X1 _0860_ ( .A1(_0201_ ), .A2(_0202_ ), .ZN(_0203_ ) );
NAND2_X1 _0861_ ( .A1(_0203_ ), .A2(_0161_ ), .ZN(_0204_ ) );
NOR2_X4 _0862_ ( .A1(_0630_ ), .A2(_0006_ ), .ZN(_0205_ ) );
OAI21_X1 _0863_ ( .A(_0200_ ), .B1(_0205_ ), .B2(_0090_ ), .ZN(_0206_ ) );
OAI21_X1 _0864_ ( .A(fanout_net_2 ), .B1(_0047_ ), .B2(_0048_ ), .ZN(_0207_ ) );
NAND2_X1 _0865_ ( .A1(_0206_ ), .A2(_0207_ ), .ZN(_0208_ ) );
NAND2_X1 _0866_ ( .A1(_0208_ ), .A2(fanout_net_4 ), .ZN(_0209_ ) );
AOI21_X1 _0867_ ( .A(_0198_ ), .B1(_0204_ ), .B2(_0209_ ), .ZN(_0210_ ) );
NOR3_X1 _0868_ ( .A1(_0098_ ), .A2(_0097_ ), .A3(_0099_ ), .ZN(_0211_ ) );
NOR3_X1 _0869_ ( .A1(_0072_ ), .A2(fanout_net_2 ), .A3(_0073_ ), .ZN(_0212_ ) );
NOR2_X1 _0870_ ( .A1(_0211_ ), .A2(_0212_ ), .ZN(_0213_ ) );
OAI211_X2 _0871_ ( .A(_0075_ ), .B(fanout_net_2 ), .C1(_0164_ ), .C2(_0078_ ), .ZN(_0214_ ) );
OAI21_X1 _0872_ ( .A(_0214_ ), .B1(_0086_ ), .B2(fanout_net_2 ), .ZN(_0215_ ) );
MUX2_X1 _0873_ ( .A(_0213_ ), .B(_0215_ ), .S(_0088_ ), .Z(_0216_ ) );
NAND2_X1 _0874_ ( .A1(_0216_ ), .A2(_0198_ ), .ZN(_0217_ ) );
AND2_X1 _0875_ ( .A1(_0069_ ), .A2(_0062_ ), .ZN(_0218_ ) );
BUF_X4 _0876_ ( .A(_0218_ ), .Z(_0219_ ) );
NAND2_X1 _0877_ ( .A1(_0217_ ), .A2(_0219_ ), .ZN(_0220_ ) );
NOR2_X1 _0878_ ( .A1(_0164_ ), .A2(_0017_ ), .ZN(_0221_ ) );
NOR3_X1 _0879_ ( .A1(_0221_ ), .A2(_0097_ ), .A3(_0612_ ), .ZN(_0222_ ) );
NOR3_X1 _0880_ ( .A1(_0052_ ), .A2(fanout_net_2 ), .A3(_0053_ ), .ZN(_0223_ ) );
NOR2_X1 _0881_ ( .A1(_0222_ ), .A2(_0223_ ), .ZN(_0224_ ) );
NAND2_X1 _0882_ ( .A1(_0224_ ), .A2(fanout_net_4 ), .ZN(_0225_ ) );
BUF_X2 _0883_ ( .A(_0060_ ), .Z(_0226_ ) );
OAI21_X1 _0884_ ( .A(_0200_ ), .B1(_0044_ ), .B2(_0045_ ), .ZN(_0227_ ) );
OAI21_X1 _0885_ ( .A(fanout_net_2 ), .B1(_0055_ ), .B2(_0056_ ), .ZN(_0228_ ) );
NAND2_X1 _0886_ ( .A1(_0227_ ), .A2(_0228_ ), .ZN(_0229_ ) );
NAND2_X1 _0887_ ( .A1(_0229_ ), .A2(_0088_ ), .ZN(_0230_ ) );
AND3_X1 _0888_ ( .A1(_0225_ ), .A2(_0226_ ), .A3(_0230_ ), .ZN(_0231_ ) );
NOR2_X1 _0889_ ( .A1(_0619_ ), .A2(_0019_ ), .ZN(_0232_ ) );
OAI21_X1 _0890_ ( .A(_0200_ ), .B1(_0232_ ), .B2(_0621_ ), .ZN(_0233_ ) );
OAI21_X1 _0891_ ( .A(fanout_net_2 ), .B1(_0631_ ), .B2(_0632_ ), .ZN(_0234_ ) );
NAND3_X1 _0892_ ( .A1(_0233_ ), .A2(_0234_ ), .A3(_0636_ ), .ZN(_0235_ ) );
NAND3_X1 _0893_ ( .A1(_0629_ ), .A2(fanout_net_4 ), .A3(_0168_ ), .ZN(_0236_ ) );
AOI21_X1 _0894_ ( .A(_0153_ ), .B1(_0235_ ), .B2(_0236_ ), .ZN(_0237_ ) );
NOR2_X1 _0895_ ( .A1(_0231_ ), .A2(_0237_ ), .ZN(_0238_ ) );
NAND2_X1 _0896_ ( .A1(_0069_ ), .A2(fanout_net_7 ), .ZN(_0239_ ) );
OAI221_X1 _0897_ ( .A(_0197_ ), .B1(_0210_ ), .B2(_0220_ ), .C1(_0238_ ), .C2(_0239_ ), .ZN(_0660_ ) );
NOR3_X1 _0898_ ( .A1(_0138_ ), .A2(_0614_ ), .A3(_0139_ ), .ZN(_0240_ ) );
NOR3_X1 _0899_ ( .A1(_0146_ ), .A2(fanout_net_2 ), .A3(_0147_ ), .ZN(_0241_ ) );
NOR2_X1 _0900_ ( .A1(_0240_ ), .A2(_0241_ ), .ZN(_0242_ ) );
NAND2_X1 _0901_ ( .A1(_0242_ ), .A2(_0625_ ), .ZN(_0243_ ) );
NOR3_X1 _0902_ ( .A1(_0118_ ), .A2(_0615_ ), .A3(_0119_ ), .ZN(_0244_ ) );
NOR3_X1 _0903_ ( .A1(_0135_ ), .A2(fanout_net_2 ), .A3(_0136_ ), .ZN(_0245_ ) );
NOR2_X1 _0904_ ( .A1(_0244_ ), .A2(_0245_ ), .ZN(_0246_ ) );
NAND2_X1 _0905_ ( .A1(_0246_ ), .A2(fanout_net_4 ), .ZN(_0247_ ) );
NAND2_X1 _0906_ ( .A1(_0243_ ), .A2(_0247_ ), .ZN(_0248_ ) );
AND2_X1 _0907_ ( .A1(_0131_ ), .A2(_0616_ ), .ZN(_0249_ ) );
INV_X1 _0908_ ( .A(_0249_ ), .ZN(_0250_ ) );
NAND2_X1 _0909_ ( .A1(_0128_ ), .A2(fanout_net_2 ), .ZN(_0251_ ) );
OAI21_X1 _0910_ ( .A(_0616_ ), .B1(_0121_ ), .B2(_0122_ ), .ZN(_0252_ ) );
NAND2_X1 _0911_ ( .A1(_0251_ ), .A2(_0252_ ), .ZN(_0253_ ) );
MUX2_X2 _0912_ ( .A(_0250_ ), .B(_0253_ ), .S(_0635_ ), .Z(_0254_ ) );
MUX2_X2 _0913_ ( .A(_0248_ ), .B(_0254_ ), .S(fanout_net_6 ), .Z(_0255_ ) );
NAND2_X1 _0914_ ( .A1(_0255_ ), .A2(fanout_net_7 ), .ZN(_0256_ ) );
INV_X1 _0915_ ( .A(_0144_ ), .ZN(_0257_ ) );
OAI211_X2 _0916_ ( .A(_0257_ ), .B(fanout_net_2 ), .C1(_0618_ ), .C2(_0009_ ), .ZN(_0258_ ) );
OAI211_X2 _0917_ ( .A(_0173_ ), .B(_0614_ ), .C1(_0618_ ), .C2(_0007_ ), .ZN(_0259_ ) );
AOI21_X1 _0918_ ( .A(_0636_ ), .B1(_0258_ ), .B2(_0259_ ), .ZN(_0260_ ) );
OAI21_X1 _0919_ ( .A(_0615_ ), .B1(_0182_ ), .B2(_0183_ ), .ZN(_0261_ ) );
NOR2_X1 _0920_ ( .A1(_0618_ ), .A2(_0005_ ), .ZN(_0262_ ) );
OAI21_X1 _0921_ ( .A(fanout_net_2 ), .B1(_0262_ ), .B2(_0175_ ), .ZN(_0263_ ) );
AND3_X1 _0922_ ( .A1(_0261_ ), .A2(_0263_ ), .A3(_0625_ ), .ZN(_0264_ ) );
OAI21_X1 _0923_ ( .A(fanout_net_6 ), .B1(_0260_ ), .B2(_0264_ ), .ZN(_0265_ ) );
NOR2_X1 _0924_ ( .A1(_0618_ ), .A2(_0030_ ), .ZN(_0266_ ) );
OAI21_X1 _0925_ ( .A(_0615_ ), .B1(_0266_ ), .B2(_0162_ ), .ZN(_0267_ ) );
OAI21_X1 _0926_ ( .A(fanout_net_3 ), .B1(_0179_ ), .B2(_0180_ ), .ZN(_0268_ ) );
NAND2_X1 _0927_ ( .A1(_0267_ ), .A2(_0268_ ), .ZN(_0269_ ) );
NAND2_X1 _0928_ ( .A1(_0269_ ), .A2(fanout_net_4 ), .ZN(_0270_ ) );
OAI211_X2 _0929_ ( .A(_0167_ ), .B(fanout_net_3 ), .C1(_0164_ ), .C2(_0028_ ), .ZN(_0271_ ) );
OAI211_X2 _0930_ ( .A(_0271_ ), .B(_0161_ ), .C1(_0159_ ), .C2(fanout_net_3 ), .ZN(_0272_ ) );
NAND3_X1 _0931_ ( .A1(_0270_ ), .A2(_0272_ ), .A3(_0106_ ), .ZN(_0273_ ) );
NAND3_X1 _0932_ ( .A1(_0265_ ), .A2(_0273_ ), .A3(_0071_ ), .ZN(_0274_ ) );
NAND3_X1 _0933_ ( .A1(_0256_ ), .A2(_0070_ ), .A3(_0274_ ), .ZN(_0275_ ) );
INV_X1 _0934_ ( .A(_0192_ ), .ZN(_0276_ ) );
BUF_X4 _0935_ ( .A(_0276_ ), .Z(_0277_ ) );
NOR2_X4 _0936_ ( .A1(_0619_ ), .A2(_0022_ ), .ZN(_0278_ ) );
NOR2_X1 _0937_ ( .A1(_0278_ ), .A2(_0158_ ), .ZN(_0279_ ) );
MUX2_X1 _0938_ ( .A(_0189_ ), .B(_0279_ ), .S(_0076_ ), .Z(_0280_ ) );
AND2_X1 _0939_ ( .A1(_0280_ ), .A2(_0161_ ), .ZN(_0281_ ) );
NAND2_X1 _0940_ ( .A1(_0281_ ), .A2(_0153_ ), .ZN(_0282_ ) );
OAI21_X1 _0941_ ( .A(_0275_ ), .B1(_0277_ ), .B2(_0282_ ), .ZN(_0663_ ) );
NAND2_X1 _0942_ ( .A1(_0050_ ), .A2(fanout_net_4 ), .ZN(_0283_ ) );
NAND3_X1 _0943_ ( .A1(_0092_ ), .A2(_0095_ ), .A3(_0624_ ), .ZN(_0284_ ) );
AND3_X1 _0944_ ( .A1(_0283_ ), .A2(fanout_net_6 ), .A3(_0284_ ), .ZN(_0285_ ) );
BUF_X4 _0945_ ( .A(_0636_ ), .Z(_0286_ ) );
AOI21_X1 _0946_ ( .A(_0286_ ), .B1(_0100_ ), .B2(_0103_ ), .ZN(_0287_ ) );
AOI21_X1 _0947_ ( .A(fanout_net_4 ), .B1(_0074_ ), .B2(_0079_ ), .ZN(_0288_ ) );
NOR3_X1 _0948_ ( .A1(_0287_ ), .A2(_0288_ ), .A3(fanout_net_6 ), .ZN(_0289_ ) );
OAI21_X1 _0949_ ( .A(_0219_ ), .B1(_0285_ ), .B2(_0289_ ), .ZN(_0290_ ) );
NAND4_X1 _0950_ ( .A1(_0168_ ), .A2(_0164_ ), .A3(fanout_net_4 ), .A4(_0000_ ), .ZN(_0291_ ) );
OR3_X4 _0951_ ( .A1(_0083_ ), .A2(_0193_ ), .A3(_0616_ ), .ZN(_0292_ ) );
NAND3_X1 _0952_ ( .A1(_0075_ ), .A2(_0130_ ), .A3(_0085_ ), .ZN(_0293_ ) );
NAND2_X1 _0953_ ( .A1(_0292_ ), .A2(_0293_ ), .ZN(_0294_ ) );
OAI21_X1 _0954_ ( .A(_0291_ ), .B1(_0294_ ), .B2(fanout_net_4 ), .ZN(_0295_ ) );
NAND3_X1 _0955_ ( .A1(_0295_ ), .A2(_0113_ ), .A3(_0192_ ), .ZN(_0296_ ) );
NAND2_X1 _0956_ ( .A1(_0058_ ), .A2(_0624_ ), .ZN(_0297_ ) );
NAND3_X1 _0957_ ( .A1(_0620_ ), .A2(_0623_ ), .A3(fanout_net_4 ), .ZN(_0298_ ) );
NAND3_X1 _0958_ ( .A1(_0297_ ), .A2(_0106_ ), .A3(_0298_ ), .ZN(_0299_ ) );
NAND3_X1 _0959_ ( .A1(_0634_ ), .A2(_0286_ ), .A3(fanout_net_6 ), .ZN(_0300_ ) );
AND2_X1 _0960_ ( .A1(_0299_ ), .A2(_0300_ ), .ZN(_0301_ ) );
OAI211_X2 _0961_ ( .A(_0290_ ), .B(_0296_ ), .C1(_0239_ ), .C2(_0301_ ), .ZN(_0664_ ) );
AND2_X1 _0962_ ( .A1(_0174_ ), .A2(_0177_ ), .ZN(_0302_ ) );
MUX2_X1 _0963_ ( .A(_0149_ ), .B(_0302_ ), .S(_0635_ ), .Z(_0303_ ) );
NAND2_X1 _0964_ ( .A1(_0303_ ), .A2(fanout_net_6 ), .ZN(_0304_ ) );
AOI21_X1 _0965_ ( .A(fanout_net_4 ), .B1(_0165_ ), .B2(_0169_ ), .ZN(_0305_ ) );
AND3_X1 _0966_ ( .A1(_0181_ ), .A2(_0184_ ), .A3(fanout_net_4 ), .ZN(_0306_ ) );
OR3_X1 _0967_ ( .A1(_0305_ ), .A2(_0306_ ), .A3(fanout_net_6 ), .ZN(_0307_ ) );
NAND3_X1 _0968_ ( .A1(_0304_ ), .A2(_0219_ ), .A3(_0307_ ), .ZN(_0308_ ) );
NAND3_X1 _0969_ ( .A1(_0189_ ), .A2(fanout_net_4 ), .A3(_0168_ ), .ZN(_0309_ ) );
OAI21_X1 _0970_ ( .A(_0130_ ), .B1(_0157_ ), .B2(_0166_ ), .ZN(_0310_ ) );
OAI21_X1 _0971_ ( .A(fanout_net_3 ), .B1(_0278_ ), .B2(_0158_ ), .ZN(_0311_ ) );
NAND2_X1 _0972_ ( .A1(_0310_ ), .A2(_0311_ ), .ZN(_0312_ ) );
OAI21_X1 _0973_ ( .A(_0309_ ), .B1(_0312_ ), .B2(fanout_net_4 ), .ZN(_0313_ ) );
NAND3_X1 _0974_ ( .A1(_0313_ ), .A2(_0113_ ), .A3(_0192_ ), .ZN(_0314_ ) );
NAND2_X1 _0975_ ( .A1(_0141_ ), .A2(_0635_ ), .ZN(_0315_ ) );
NAND2_X1 _0976_ ( .A1(_0124_ ), .A2(fanout_net_4 ), .ZN(_0316_ ) );
BUF_X2 _0977_ ( .A(_0060_ ), .Z(_0317_ ) );
AND3_X1 _0978_ ( .A1(_0315_ ), .A2(_0316_ ), .A3(_0317_ ), .ZN(_0318_ ) );
NOR3_X1 _0979_ ( .A1(_0132_ ), .A2(fanout_net_4 ), .A3(_0226_ ), .ZN(_0319_ ) );
NOR2_X1 _0980_ ( .A1(_0318_ ), .A2(_0319_ ), .ZN(_0320_ ) );
OAI211_X2 _0981_ ( .A(_0308_ ), .B(_0314_ ), .C1(_0239_ ), .C2(_0320_ ), .ZN(_0665_ ) );
NAND2_X1 _0982_ ( .A1(_0194_ ), .A2(_0195_ ), .ZN(_0321_ ) );
NAND2_X1 _0983_ ( .A1(_0321_ ), .A2(fanout_net_4 ), .ZN(_0322_ ) );
NOR2_X1 _0984_ ( .A1(_0077_ ), .A2(_0027_ ), .ZN(_0323_ ) );
OAI21_X1 _0985_ ( .A(_0097_ ), .B1(_0323_ ), .B2(_0073_ ), .ZN(_0324_ ) );
NAND3_X1 _0986_ ( .A1(_0075_ ), .A2(fanout_net_3 ), .A3(_0085_ ), .ZN(_0325_ ) );
NAND2_X1 _0987_ ( .A1(_0324_ ), .A2(_0325_ ), .ZN(_0326_ ) );
OAI21_X1 _0988_ ( .A(_0322_ ), .B1(fanout_net_4 ), .B2(_0326_ ), .ZN(_0327_ ) );
NAND3_X1 _0989_ ( .A1(_0327_ ), .A2(_0113_ ), .A3(_0192_ ), .ZN(_0328_ ) );
NAND2_X1 _0990_ ( .A1(_0224_ ), .A2(_0161_ ), .ZN(_0329_ ) );
NAND2_X1 _0991_ ( .A1(_0233_ ), .A2(_0234_ ), .ZN(_0330_ ) );
NAND2_X1 _0992_ ( .A1(_0330_ ), .A2(fanout_net_4 ), .ZN(_0331_ ) );
NAND3_X1 _0993_ ( .A1(_0329_ ), .A2(_0331_ ), .A3(_0226_ ), .ZN(_0332_ ) );
NAND4_X1 _0994_ ( .A1(_0629_ ), .A2(_0286_ ), .A3(_0168_ ), .A4(fanout_net_6 ), .ZN(_0333_ ) );
AND2_X1 _0995_ ( .A1(_0332_ ), .A2(_0333_ ), .ZN(_0334_ ) );
MUX2_X1 _0996_ ( .A(_0203_ ), .B(_0213_ ), .S(_0161_ ), .Z(_0335_ ) );
NAND2_X1 _0997_ ( .A1(_0335_ ), .A2(_0198_ ), .ZN(_0336_ ) );
NAND2_X1 _0998_ ( .A1(_0336_ ), .A2(_0219_ ), .ZN(_0337_ ) );
NAND2_X1 _0999_ ( .A1(_0208_ ), .A2(_0088_ ), .ZN(_0338_ ) );
NAND2_X1 _1000_ ( .A1(_0229_ ), .A2(fanout_net_4 ), .ZN(_0339_ ) );
AOI21_X1 _1001_ ( .A(_0198_ ), .B1(_0338_ ), .B2(_0339_ ), .ZN(_0340_ ) );
OAI221_X1 _1002_ ( .A(_0328_ ), .B1(_0334_ ), .B2(_0239_ ), .C1(_0337_ ), .C2(_0340_ ), .ZN(_0666_ ) );
INV_X1 _1003_ ( .A(_0069_ ), .ZN(_0341_ ) );
NAND2_X1 _1004_ ( .A1(_0242_ ), .A2(fanout_net_4 ), .ZN(_0342_ ) );
NAND3_X1 _1005_ ( .A1(_0258_ ), .A2(_0259_ ), .A3(_0624_ ), .ZN(_0343_ ) );
AND3_X2 _1006_ ( .A1(_0342_ ), .A2(fanout_net_6 ), .A3(_0343_ ), .ZN(_0344_ ) );
NAND3_X1 _1007_ ( .A1(_0261_ ), .A2(_0263_ ), .A3(fanout_net_5 ), .ZN(_0345_ ) );
OAI21_X1 _1008_ ( .A(_0345_ ), .B1(_0269_ ), .B2(fanout_net_5 ), .ZN(_0346_ ) );
AOI211_X2 _1009_ ( .A(fanout_net_7 ), .B(_0344_ ), .C1(_0041_ ), .C2(_0346_ ), .ZN(_0347_ ) );
NAND2_X1 _1010_ ( .A1(_0253_ ), .A2(fanout_net_5 ), .ZN(_0348_ ) );
NAND2_X1 _1011_ ( .A1(_0246_ ), .A2(_0624_ ), .ZN(_0349_ ) );
NAND3_X1 _1012_ ( .A1(_0348_ ), .A2(_0041_ ), .A3(_0349_ ), .ZN(_0350_ ) );
NAND4_X1 _1013_ ( .A1(_0131_ ), .A2(_0635_ ), .A3(_0097_ ), .A4(fanout_net_6 ), .ZN(_0351_ ) );
AND2_X1 _1014_ ( .A1(_0350_ ), .A2(_0351_ ), .ZN(_0352_ ) );
AOI211_X2 _1015_ ( .A(_0341_ ), .B(_0347_ ), .C1(fanout_net_7 ), .C2(_0352_ ), .ZN(_0353_ ) );
OAI211_X2 _1016_ ( .A(_0163_ ), .B(_0130_ ), .C1(_0164_ ), .C2(_0028_ ), .ZN(_0354_ ) );
OAI211_X2 _1017_ ( .A(_0167_ ), .B(fanout_net_3 ), .C1(_0164_ ), .C2(_0026_ ), .ZN(_0355_ ) );
NAND2_X1 _1018_ ( .A1(_0354_ ), .A2(_0355_ ), .ZN(_0356_ ) );
MUX2_X2 _1019_ ( .A(_0356_ ), .B(_0280_ ), .S(fanout_net_5 ), .Z(_0357_ ) );
AND3_X1 _1020_ ( .A1(_0357_ ), .A2(_0198_ ), .A3(_0192_ ), .ZN(_0358_ ) );
OR2_X1 _1021_ ( .A1(_0353_ ), .A2(_0358_ ), .ZN(_0667_ ) );
AND3_X1 _1022_ ( .A1(_0051_ ), .A2(_0059_ ), .A3(fanout_net_6 ), .ZN(_0359_ ) );
AOI21_X1 _1023_ ( .A(_0359_ ), .B1(_0106_ ), .B2(_0105_ ), .ZN(_0360_ ) );
AOI21_X1 _1024_ ( .A(_0341_ ), .B1(_0360_ ), .B2(_0071_ ), .ZN(_0361_ ) );
NOR2_X1 _1025_ ( .A1(_0637_ ), .A2(fanout_net_6 ), .ZN(_0362_ ) );
OAI21_X1 _1026_ ( .A(_0361_ ), .B1(_0071_ ), .B2(_0362_ ), .ZN(_0363_ ) );
INV_X1 _1027_ ( .A(_0116_ ), .ZN(_0364_ ) );
NAND2_X1 _1028_ ( .A1(_0294_ ), .A2(fanout_net_5 ), .ZN(_0365_ ) );
OAI21_X1 _1029_ ( .A(_0130_ ), .B1(_0072_ ), .B2(_0099_ ), .ZN(_0366_ ) );
OAI21_X1 _1030_ ( .A(fanout_net_3 ), .B1(_0323_ ), .B2(_0073_ ), .ZN(_0367_ ) );
NAND2_X1 _1031_ ( .A1(_0366_ ), .A2(_0367_ ), .ZN(_0368_ ) );
NAND2_X1 _1032_ ( .A1(_0368_ ), .A2(_0625_ ), .ZN(_0369_ ) );
NAND2_X1 _1033_ ( .A1(_0365_ ), .A2(_0369_ ), .ZN(_0370_ ) );
MUX2_X2 _1034_ ( .A(_0364_ ), .B(_0370_ ), .S(_0042_ ), .Z(_0371_ ) );
OAI21_X1 _1035_ ( .A(_0363_ ), .B1(_0277_ ), .B2(_0371_ ), .ZN(_0668_ ) );
NOR3_X1 _1036_ ( .A1(_0133_ ), .A2(fanout_net_6 ), .A3(_0063_ ), .ZN(_0372_ ) );
NAND3_X1 _1037_ ( .A1(_0142_ ), .A2(fanout_net_6 ), .A3(_0150_ ), .ZN(_0373_ ) );
OAI21_X1 _1038_ ( .A(_0226_ ), .B1(_0178_ ), .B2(_0185_ ), .ZN(_0374_ ) );
AOI21_X1 _1039_ ( .A(fanout_net_7 ), .B1(_0373_ ), .B2(_0374_ ), .ZN(_0375_ ) );
OAI21_X1 _1040_ ( .A(_0070_ ), .B1(_0372_ ), .B2(_0375_ ), .ZN(_0376_ ) );
NOR2_X1 _1041_ ( .A1(_0077_ ), .A2(_0028_ ), .ZN(_0377_ ) );
NOR3_X1 _1042_ ( .A1(_0377_ ), .A2(_0076_ ), .A3(_0162_ ), .ZN(_0378_ ) );
NOR3_X1 _1043_ ( .A1(_0266_ ), .A2(fanout_net_3 ), .A3(_0180_ ), .ZN(_0379_ ) );
NOR2_X1 _1044_ ( .A1(_0378_ ), .A2(_0379_ ), .ZN(_0380_ ) );
NAND2_X1 _1045_ ( .A1(_0380_ ), .A2(_0625_ ), .ZN(_0381_ ) );
NAND2_X1 _1046_ ( .A1(_0312_ ), .A2(fanout_net_5 ), .ZN(_0382_ ) );
NAND3_X1 _1047_ ( .A1(_0381_ ), .A2(_0382_ ), .A3(_0317_ ), .ZN(_0383_ ) );
NAND4_X1 _1048_ ( .A1(_0189_ ), .A2(_0286_ ), .A3(_0168_ ), .A4(fanout_net_6 ), .ZN(_0384_ ) );
AND2_X1 _1049_ ( .A1(_0383_ ), .A2(_0384_ ), .ZN(_0385_ ) );
OAI21_X1 _1050_ ( .A(_0376_ ), .B1(_0277_ ), .B2(_0385_ ), .ZN(_0669_ ) );
AOI21_X1 _1051_ ( .A(fanout_net_6 ), .B1(_0204_ ), .B2(_0209_ ), .ZN(_0386_ ) );
AOI21_X1 _1052_ ( .A(_0317_ ), .B1(_0225_ ), .B2(_0230_ ), .ZN(_0387_ ) );
NOR3_X1 _1053_ ( .A1(_0386_ ), .A2(_0387_ ), .A3(fanout_net_7 ), .ZN(_0388_ ) );
AOI211_X4 _1054_ ( .A(fanout_net_6 ), .B(_0063_ ), .C1(_0235_ ), .C2(_0236_ ), .ZN(_0389_ ) );
OAI21_X1 _1055_ ( .A(_0070_ ), .B1(_0388_ ), .B2(_0389_ ), .ZN(_0390_ ) );
NOR3_X1 _1056_ ( .A1(_0072_ ), .A2(_0200_ ), .A3(_0099_ ), .ZN(_0391_ ) );
NOR3_X1 _1057_ ( .A1(_0098_ ), .A2(fanout_net_3 ), .A3(_0102_ ), .ZN(_0392_ ) );
NOR2_X1 _1058_ ( .A1(_0391_ ), .A2(_0392_ ), .ZN(_0393_ ) );
NAND2_X1 _1059_ ( .A1(_0393_ ), .A2(_0161_ ), .ZN(_0394_ ) );
NAND2_X1 _1060_ ( .A1(_0326_ ), .A2(fanout_net_5 ), .ZN(_0395_ ) );
NAND3_X1 _1061_ ( .A1(_0394_ ), .A2(_0395_ ), .A3(_0226_ ), .ZN(_0396_ ) );
NAND3_X1 _1062_ ( .A1(_0321_ ), .A2(_0286_ ), .A3(fanout_net_6 ), .ZN(_0397_ ) );
AND2_X1 _1063_ ( .A1(_0396_ ), .A2(_0397_ ), .ZN(_0398_ ) );
OAI21_X1 _1064_ ( .A(_0390_ ), .B1(_0277_ ), .B2(_0398_ ), .ZN(_0639_ ) );
NOR3_X1 _1065_ ( .A1(_0254_ ), .A2(fanout_net_6 ), .A3(_0063_ ), .ZN(_0399_ ) );
AOI21_X1 _1066_ ( .A(_0317_ ), .B1(_0243_ ), .B2(_0247_ ), .ZN(_0400_ ) );
NOR3_X1 _1067_ ( .A1(_0260_ ), .A2(_0264_ ), .A3(fanout_net_6 ), .ZN(_0401_ ) );
NOR3_X1 _1068_ ( .A1(_0400_ ), .A2(_0401_ ), .A3(fanout_net_7 ), .ZN(_0402_ ) );
OAI21_X1 _1069_ ( .A(_0070_ ), .B1(_0399_ ), .B2(_0402_ ), .ZN(_0403_ ) );
NAND3_X1 _1070_ ( .A1(_0280_ ), .A2(_0286_ ), .A3(fanout_net_6 ), .ZN(_0404_ ) );
OAI21_X1 _1071_ ( .A(_0130_ ), .B1(_0179_ ), .B2(_0183_ ), .ZN(_0405_ ) );
OAI21_X1 _1072_ ( .A(fanout_net_3 ), .B1(_0266_ ), .B2(_0180_ ), .ZN(_0406_ ) );
NAND2_X1 _1073_ ( .A1(_0405_ ), .A2(_0406_ ), .ZN(_0407_ ) );
NAND2_X1 _1074_ ( .A1(_0407_ ), .A2(_0625_ ), .ZN(_0408_ ) );
NAND3_X1 _1075_ ( .A1(_0354_ ), .A2(_0355_ ), .A3(fanout_net_5 ), .ZN(_0409_ ) );
NAND3_X1 _1076_ ( .A1(_0408_ ), .A2(_0226_ ), .A3(_0409_ ), .ZN(_0410_ ) );
AND2_X1 _1077_ ( .A1(_0404_ ), .A2(_0410_ ), .ZN(_0411_ ) );
OAI21_X1 _1078_ ( .A(_0403_ ), .B1(_0277_ ), .B2(_0411_ ), .ZN(_0640_ ) );
NAND3_X1 _1079_ ( .A1(_0283_ ), .A2(_0041_ ), .A3(_0284_ ), .ZN(_0412_ ) );
NAND3_X1 _1080_ ( .A1(_0297_ ), .A2(fanout_net_6 ), .A3(_0298_ ), .ZN(_0413_ ) );
AND3_X1 _1081_ ( .A1(_0412_ ), .A2(_0413_ ), .A3(_0063_ ), .ZN(_0414_ ) );
AND2_X1 _1082_ ( .A1(_0634_ ), .A2(_0635_ ), .ZN(_0415_ ) );
NAND2_X1 _1083_ ( .A1(_0415_ ), .A2(_0060_ ), .ZN(_0416_ ) );
AOI211_X2 _1084_ ( .A(_0341_ ), .B(_0414_ ), .C1(fanout_net_7 ), .C2(_0416_ ), .ZN(_0417_ ) );
NOR3_X1 _1085_ ( .A1(_0098_ ), .A2(_0616_ ), .A3(_0102_ ), .ZN(_0418_ ) );
NOR3_X1 _1086_ ( .A1(_0101_ ), .A2(fanout_net_3 ), .A3(_0093_ ), .ZN(_0419_ ) );
OR3_X1 _1087_ ( .A1(_0418_ ), .A2(_0419_ ), .A3(fanout_net_5 ), .ZN(_0420_ ) );
NAND2_X1 _1088_ ( .A1(_0368_ ), .A2(fanout_net_5 ), .ZN(_0421_ ) );
NAND2_X2 _1089_ ( .A1(_0420_ ), .A2(_0421_ ), .ZN(_0422_ ) );
NAND2_X1 _1090_ ( .A1(_0422_ ), .A2(_0042_ ), .ZN(_0423_ ) );
OAI21_X1 _1091_ ( .A(_0423_ ), .B1(_0106_ ), .B2(_0295_ ), .ZN(_0424_ ) );
NOR2_X1 _1092_ ( .A1(_0424_ ), .A2(_0276_ ), .ZN(_0425_ ) );
OR2_X1 _1093_ ( .A1(_0417_ ), .A2(_0425_ ), .ZN(_0641_ ) );
AOI21_X1 _1094_ ( .A(_0060_ ), .B1(_0315_ ), .B2(_0316_ ), .ZN(_0426_ ) );
AOI211_X2 _1095_ ( .A(fanout_net_7 ), .B(_0426_ ), .C1(_0042_ ), .C2(_0303_ ), .ZN(_0427_ ) );
NOR4_X1 _1096_ ( .A1(_0132_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .A4(_0063_ ), .ZN(_0428_ ) );
OAI21_X1 _1097_ ( .A(_0070_ ), .B1(_0427_ ), .B2(_0428_ ), .ZN(_0429_ ) );
NAND2_X1 _1098_ ( .A1(_0380_ ), .A2(fanout_net_5 ), .ZN(_0430_ ) );
OAI21_X1 _1099_ ( .A(_0130_ ), .B1(_0182_ ), .B2(_0175_ ), .ZN(_0431_ ) );
OAI21_X1 _1100_ ( .A(fanout_net_3 ), .B1(_0179_ ), .B2(_0183_ ), .ZN(_0432_ ) );
NAND2_X1 _1101_ ( .A1(_0431_ ), .A2(_0432_ ), .ZN(_0433_ ) );
NAND2_X1 _1102_ ( .A1(_0433_ ), .A2(_0636_ ), .ZN(_0434_ ) );
NAND2_X1 _1103_ ( .A1(_0430_ ), .A2(_0434_ ), .ZN(_0435_ ) );
NAND2_X1 _1104_ ( .A1(_0435_ ), .A2(_0226_ ), .ZN(_0436_ ) );
OAI21_X1 _1105_ ( .A(_0436_ ), .B1(_0313_ ), .B2(_0153_ ), .ZN(_0437_ ) );
OAI21_X1 _1106_ ( .A(_0429_ ), .B1(_0277_ ), .B2(_0437_ ), .ZN(_0642_ ) );
AOI21_X1 _1107_ ( .A(_0226_ ), .B1(_0329_ ), .B2(_0331_ ), .ZN(_0438_ ) );
AOI21_X1 _1108_ ( .A(fanout_net_6 ), .B1(_0338_ ), .B2(_0339_ ), .ZN(_0439_ ) );
NOR3_X1 _1109_ ( .A1(_0438_ ), .A2(_0439_ ), .A3(fanout_net_7 ), .ZN(_0440_ ) );
AND3_X1 _1110_ ( .A1(_0629_ ), .A2(_0636_ ), .A3(_0168_ ), .ZN(_0441_ ) );
AND3_X1 _1111_ ( .A1(_0441_ ), .A2(_0106_ ), .A3(fanout_net_7 ), .ZN(_0442_ ) );
OAI21_X1 _1112_ ( .A(_0070_ ), .B1(_0440_ ), .B2(_0442_ ), .ZN(_0443_ ) );
NAND2_X1 _1113_ ( .A1(_0327_ ), .A2(fanout_net_6 ), .ZN(_0444_ ) );
NAND2_X1 _1114_ ( .A1(_0393_ ), .A2(fanout_net_5 ), .ZN(_0445_ ) );
OAI21_X1 _1115_ ( .A(_0200_ ), .B1(_0199_ ), .B2(_0090_ ), .ZN(_0446_ ) );
OAI21_X1 _1116_ ( .A(fanout_net_3 ), .B1(_0101_ ), .B2(_0093_ ), .ZN(_0447_ ) );
NAND2_X1 _1117_ ( .A1(_0446_ ), .A2(_0447_ ), .ZN(_0448_ ) );
NAND2_X1 _1118_ ( .A1(_0448_ ), .A2(_0161_ ), .ZN(_0449_ ) );
NAND3_X1 _1119_ ( .A1(_0445_ ), .A2(_0153_ ), .A3(_0449_ ), .ZN(_0450_ ) );
AND2_X1 _1120_ ( .A1(_0444_ ), .A2(_0450_ ), .ZN(_0451_ ) );
OAI21_X1 _1121_ ( .A(_0443_ ), .B1(_0451_ ), .B2(_0277_ ), .ZN(_0643_ ) );
AOI21_X1 _1122_ ( .A(_0317_ ), .B1(_0348_ ), .B2(_0349_ ), .ZN(_0452_ ) );
AOI21_X1 _1123_ ( .A(fanout_net_6 ), .B1(_0342_ ), .B2(_0343_ ), .ZN(_0453_ ) );
NOR3_X1 _1124_ ( .A1(_0452_ ), .A2(_0453_ ), .A3(fanout_net_7 ), .ZN(_0454_ ) );
AND3_X1 _1125_ ( .A1(_0131_ ), .A2(_0088_ ), .A3(_0168_ ), .ZN(_0455_ ) );
AND3_X1 _1126_ ( .A1(_0455_ ), .A2(_0106_ ), .A3(fanout_net_7 ), .ZN(_0456_ ) );
OAI21_X1 _1127_ ( .A(_0070_ ), .B1(_0454_ ), .B2(_0456_ ), .ZN(_0457_ ) );
NAND2_X1 _1128_ ( .A1(_0357_ ), .A2(fanout_net_6 ), .ZN(_0458_ ) );
NOR3_X1 _1129_ ( .A1(_0182_ ), .A2(_0076_ ), .A3(_0175_ ), .ZN(_0459_ ) );
NOR3_X1 _1130_ ( .A1(_0262_ ), .A2(fanout_net_3 ), .A3(_0172_ ), .ZN(_0460_ ) );
NOR2_X1 _1131_ ( .A1(_0459_ ), .A2(_0460_ ), .ZN(_0461_ ) );
NAND2_X1 _1132_ ( .A1(_0461_ ), .A2(_0161_ ), .ZN(_0462_ ) );
NAND2_X1 _1133_ ( .A1(_0407_ ), .A2(fanout_net_5 ), .ZN(_0463_ ) );
NAND3_X1 _1134_ ( .A1(_0462_ ), .A2(_0463_ ), .A3(_0226_ ), .ZN(_0464_ ) );
AND2_X2 _1135_ ( .A1(_0458_ ), .A2(_0464_ ), .ZN(_0465_ ) );
OAI21_X1 _1136_ ( .A(_0457_ ), .B1(_0465_ ), .B2(_0277_ ), .ZN(_0644_ ) );
OAI21_X2 _1137_ ( .A(fanout_net_5 ), .B1(_0418_ ), .B2(_0419_ ), .ZN(_0466_ ) );
NOR3_X1 _1138_ ( .A1(_0199_ ), .A2(_0616_ ), .A3(_0090_ ), .ZN(_0467_ ) );
NOR3_X1 _1139_ ( .A1(_0205_ ), .A2(fanout_net_3 ), .A3(_0048_ ), .ZN(_0468_ ) );
OAI21_X1 _1140_ ( .A(_0635_ ), .B1(_0467_ ), .B2(_0468_ ), .ZN(_0469_ ) );
AND3_X1 _1141_ ( .A1(_0466_ ), .A2(_0469_ ), .A3(_0060_ ), .ZN(_0470_ ) );
AOI211_X2 _1142_ ( .A(fanout_net_7 ), .B(_0470_ ), .C1(_0035_ ), .C2(_0370_ ), .ZN(_0471_ ) );
AND3_X1 _1143_ ( .A1(_0116_ ), .A2(_0153_ ), .A3(fanout_net_7 ), .ZN(_0472_ ) );
OAI21_X1 _1144_ ( .A(_0112_ ), .B1(_0471_ ), .B2(_0472_ ), .ZN(_0473_ ) );
OAI21_X1 _1145_ ( .A(_0219_ ), .B1(_0043_ ), .B2(_0061_ ), .ZN(_0474_ ) );
NAND2_X1 _1146_ ( .A1(_0473_ ), .A2(_0474_ ), .ZN(_0645_ ) );
AOI21_X1 _1147_ ( .A(_0060_ ), .B1(_0381_ ), .B2(_0382_ ), .ZN(_0475_ ) );
OAI211_X2 _1148_ ( .A(_0173_ ), .B(fanout_net_3 ), .C1(_0077_ ), .C2(_0005_ ), .ZN(_0476_ ) );
OAI211_X2 _1149_ ( .A(_0257_ ), .B(_0616_ ), .C1(_0077_ ), .C2(_0007_ ), .ZN(_0477_ ) );
AND2_X1 _1150_ ( .A1(_0476_ ), .A2(_0477_ ), .ZN(_0478_ ) );
MUX2_X1 _1151_ ( .A(_0433_ ), .B(_0478_ ), .S(_0635_ ), .Z(_0479_ ) );
AOI211_X2 _1152_ ( .A(fanout_net_7 ), .B(_0475_ ), .C1(_0317_ ), .C2(_0479_ ), .ZN(_0480_ ) );
AND3_X1 _1153_ ( .A1(_0190_ ), .A2(_0153_ ), .A3(fanout_net_7 ), .ZN(_0481_ ) );
OAI21_X1 _1154_ ( .A(_0112_ ), .B1(_0480_ ), .B2(_0481_ ), .ZN(_0482_ ) );
OAI21_X1 _1155_ ( .A(_0219_ ), .B1(_0134_ ), .B2(_0151_ ), .ZN(_0483_ ) );
NAND2_X1 _1156_ ( .A1(_0482_ ), .A2(_0483_ ), .ZN(_0646_ ) );
AOI21_X1 _1157_ ( .A(_0317_ ), .B1(_0394_ ), .B2(_0395_ ), .ZN(_0484_ ) );
OAI21_X1 _1158_ ( .A(_0200_ ), .B1(_0047_ ), .B2(_0045_ ), .ZN(_0485_ ) );
OAI21_X1 _1159_ ( .A(fanout_net_3 ), .B1(_0205_ ), .B2(_0048_ ), .ZN(_0486_ ) );
NAND2_X1 _1160_ ( .A1(_0485_ ), .A2(_0486_ ), .ZN(_0487_ ) );
NAND2_X1 _1161_ ( .A1(_0487_ ), .A2(_0088_ ), .ZN(_0488_ ) );
NAND2_X1 _1162_ ( .A1(_0448_ ), .A2(fanout_net_5 ), .ZN(_0489_ ) );
AOI21_X1 _1163_ ( .A(_0035_ ), .B1(_0488_ ), .B2(_0489_ ), .ZN(_0490_ ) );
NOR3_X1 _1164_ ( .A1(_0484_ ), .A2(_0490_ ), .A3(fanout_net_7 ), .ZN(_0491_ ) );
AND4_X1 _1165_ ( .A1(_0286_ ), .A2(_0321_ ), .A3(_0317_ ), .A4(fanout_net_7 ), .ZN(_0492_ ) );
OAI21_X1 _1166_ ( .A(_0112_ ), .B1(_0491_ ), .B2(_0492_ ), .ZN(_0493_ ) );
INV_X2 _1167_ ( .A(_0219_ ), .ZN(_0494_ ) );
OAI21_X1 _1168_ ( .A(_0493_ ), .B1(_0494_ ), .B2(_0238_ ), .ZN(_0647_ ) );
NAND3_X1 _1169_ ( .A1(_0408_ ), .A2(_0035_ ), .A3(_0409_ ), .ZN(_0495_ ) );
NOR2_X4 _1170_ ( .A1(_0077_ ), .A2(_0007_ ), .ZN(_0496_ ) );
NOR3_X4 _1171_ ( .A1(_0496_ ), .A2(_0076_ ), .A3(_0144_ ), .ZN(_0497_ ) );
NOR3_X1 _1172_ ( .A1(_0143_ ), .A2(fanout_net_3 ), .A3(_0147_ ), .ZN(_0498_ ) );
NOR2_X1 _1173_ ( .A1(_0497_ ), .A2(_0498_ ), .ZN(_0499_ ) );
MUX2_X2 _1174_ ( .A(_0499_ ), .B(_0461_ ), .S(fanout_net_5 ), .Z(_0500_ ) );
OAI21_X1 _1175_ ( .A(_0495_ ), .B1(_0500_ ), .B2(_0035_ ), .ZN(_0501_ ) );
OAI21_X1 _1176_ ( .A(_0111_ ), .B1(_0501_ ), .B2(fanout_net_7 ), .ZN(_0502_ ) );
AOI21_X1 _1177_ ( .A(_0502_ ), .B1(fanout_net_7 ), .B2(_0282_ ), .ZN(_0503_ ) );
NOR2_X1 _1178_ ( .A1(_0255_ ), .A2(_0494_ ), .ZN(_0504_ ) );
OR2_X1 _1179_ ( .A1(_0503_ ), .A2(_0504_ ), .ZN(_0648_ ) );
OR3_X4 _1180_ ( .A1(_0047_ ), .A2(_0614_ ), .A3(_0045_ ), .ZN(_0505_ ) );
OR3_X2 _1181_ ( .A1(_0044_ ), .A2(fanout_net_3 ), .A3(_0056_ ), .ZN(_0506_ ) );
AND2_X2 _1182_ ( .A1(_0505_ ), .A2(_0506_ ), .ZN(_0507_ ) );
OR2_X4 _1183_ ( .A1(_0507_ ), .A2(fanout_net_5 ), .ZN(_0508_ ) );
OAI21_X1 _1184_ ( .A(fanout_net_5 ), .B1(_0467_ ), .B2(_0468_ ), .ZN(_0509_ ) );
AND3_X2 _1185_ ( .A1(_0508_ ), .A2(_0041_ ), .A3(_0509_ ), .ZN(_0510_ ) );
AOI211_X2 _1186_ ( .A(fanout_net_7 ), .B(_0510_ ), .C1(_0035_ ), .C2(_0422_ ), .ZN(_0511_ ) );
AND3_X1 _1187_ ( .A1(_0295_ ), .A2(_0106_ ), .A3(fanout_net_7 ), .ZN(_0512_ ) );
OAI21_X1 _1188_ ( .A(_0112_ ), .B1(_0511_ ), .B2(_0512_ ), .ZN(_0513_ ) );
OAI21_X1 _1189_ ( .A(_0513_ ), .B1(_0494_ ), .B2(_0301_ ), .ZN(_0650_ ) );
AND2_X1 _1190_ ( .A1(_0313_ ), .A2(_0317_ ), .ZN(_0514_ ) );
OAI21_X1 _1191_ ( .A(_0063_ ), .B1(_0435_ ), .B2(_0198_ ), .ZN(_0515_ ) );
AND3_X1 _1192_ ( .A1(_0476_ ), .A2(_0477_ ), .A3(fanout_net_5 ), .ZN(_0516_ ) );
OAI21_X1 _1193_ ( .A(_0097_ ), .B1(_0146_ ), .B2(_0139_ ), .ZN(_0517_ ) );
OAI21_X1 _1194_ ( .A(fanout_net_3 ), .B1(_0143_ ), .B2(_0147_ ), .ZN(_0518_ ) );
AOI21_X1 _1195_ ( .A(fanout_net_5 ), .B1(_0517_ ), .B2(_0518_ ), .ZN(_0519_ ) );
NOR3_X1 _1196_ ( .A1(_0516_ ), .A2(_0035_ ), .A3(_0519_ ), .ZN(_0520_ ) );
OAI221_X1 _1197_ ( .A(_0111_ ), .B1(_0071_ ), .B2(_0514_ ), .C1(_0515_ ), .C2(_0520_ ), .ZN(_0521_ ) );
OAI21_X1 _1198_ ( .A(_0521_ ), .B1(_0494_ ), .B2(_0320_ ), .ZN(_0651_ ) );
AOI21_X1 _1199_ ( .A(_0317_ ), .B1(_0445_ ), .B2(_0449_ ), .ZN(_0522_ ) );
OAI21_X1 _1200_ ( .A(_0200_ ), .B1(_0055_ ), .B2(_0053_ ), .ZN(_0523_ ) );
OAI21_X1 _1201_ ( .A(fanout_net_3 ), .B1(_0044_ ), .B2(_0056_ ), .ZN(_0524_ ) );
NAND2_X1 _1202_ ( .A1(_0523_ ), .A2(_0524_ ), .ZN(_0525_ ) );
NAND2_X1 _1203_ ( .A1(_0525_ ), .A2(_0088_ ), .ZN(_0526_ ) );
NAND2_X1 _1204_ ( .A1(_0487_ ), .A2(fanout_net_5 ), .ZN(_0527_ ) );
AOI21_X1 _1205_ ( .A(_0035_ ), .B1(_0526_ ), .B2(_0527_ ), .ZN(_0528_ ) );
NOR3_X1 _1206_ ( .A1(_0522_ ), .A2(_0528_ ), .A3(fanout_net_7 ), .ZN(_0529_ ) );
AND3_X1 _1207_ ( .A1(_0327_ ), .A2(_0106_ ), .A3(fanout_net_7 ), .ZN(_0530_ ) );
OAI21_X1 _1208_ ( .A(_0112_ ), .B1(_0529_ ), .B2(_0530_ ), .ZN(_0531_ ) );
OAI21_X1 _1209_ ( .A(_0531_ ), .B1(_0494_ ), .B2(_0334_ ), .ZN(_0652_ ) );
AND3_X1 _1210_ ( .A1(_0357_ ), .A2(_0153_ ), .A3(fanout_net_7 ), .ZN(_0532_ ) );
NAND2_X1 _1211_ ( .A1(_0499_ ), .A2(fanout_net_5 ), .ZN(_0533_ ) );
OAI21_X1 _1212_ ( .A(_0200_ ), .B1(_0138_ ), .B2(_0136_ ), .ZN(_0534_ ) );
OAI21_X1 _1213_ ( .A(fanout_net_3 ), .B1(_0146_ ), .B2(_0139_ ), .ZN(_0535_ ) );
NAND2_X1 _1214_ ( .A1(_0534_ ), .A2(_0535_ ), .ZN(_0536_ ) );
NAND2_X1 _1215_ ( .A1(_0536_ ), .A2(_0161_ ), .ZN(_0537_ ) );
NAND3_X1 _1216_ ( .A1(_0533_ ), .A2(_0226_ ), .A3(_0537_ ), .ZN(_0538_ ) );
NAND3_X1 _1217_ ( .A1(_0462_ ), .A2(_0463_ ), .A3(_0035_ ), .ZN(_0539_ ) );
AOI21_X1 _1218_ ( .A(fanout_net_7 ), .B1(_0538_ ), .B2(_0539_ ), .ZN(_0540_ ) );
OAI21_X1 _1219_ ( .A(_0112_ ), .B1(_0532_ ), .B2(_0540_ ), .ZN(_0541_ ) );
OAI21_X1 _1220_ ( .A(_0541_ ), .B1(_0494_ ), .B2(_0352_ ), .ZN(_0653_ ) );
OR3_X4 _1221_ ( .A1(_0055_ ), .A2(_0615_ ), .A3(_0053_ ), .ZN(_0542_ ) );
NOR2_X2 _1222_ ( .A1(_0052_ ), .A2(_0612_ ), .ZN(_0543_ ) );
INV_X2 _1223_ ( .A(_0543_ ), .ZN(_0544_ ) );
OAI211_X2 _1224_ ( .A(_0542_ ), .B(_0624_ ), .C1(_0544_ ), .C2(fanout_net_3 ), .ZN(_0545_ ) );
NAND3_X1 _1225_ ( .A1(_0505_ ), .A2(_0506_ ), .A3(fanout_net_5 ), .ZN(_0546_ ) );
AND3_X1 _1226_ ( .A1(_0545_ ), .A2(_0041_ ), .A3(_0546_ ), .ZN(_0547_ ) );
AOI21_X1 _1227_ ( .A(_0041_ ), .B1(_0466_ ), .B2(_0469_ ), .ZN(_0548_ ) );
OR3_X2 _1228_ ( .A1(_0547_ ), .A2(fanout_net_7 ), .A3(_0548_ ), .ZN(_0549_ ) );
NAND2_X1 _1229_ ( .A1(_0549_ ), .A2(_0111_ ), .ZN(_0550_ ) );
AOI21_X1 _1230_ ( .A(_0550_ ), .B1(fanout_net_7 ), .B2(_0371_ ), .ZN(_0551_ ) );
NOR3_X1 _1231_ ( .A1(_0637_ ), .A2(_0035_ ), .A3(_0494_ ), .ZN(_0552_ ) );
OR2_X1 _1232_ ( .A1(_0551_ ), .A2(_0552_ ), .ZN(_0654_ ) );
OR3_X1 _1233_ ( .A1(_0138_ ), .A2(_0076_ ), .A3(_0136_ ), .ZN(_0553_ ) );
OR3_X1 _1234_ ( .A1(_0135_ ), .A2(fanout_net_3 ), .A3(_0119_ ), .ZN(_0554_ ) );
AND3_X1 _1235_ ( .A1(_0553_ ), .A2(_0554_ ), .A3(_0625_ ), .ZN(_0555_ ) );
AOI21_X1 _1236_ ( .A(_0636_ ), .B1(_0517_ ), .B2(_0518_ ), .ZN(_0556_ ) );
OAI21_X1 _1237_ ( .A(_0042_ ), .B1(_0555_ ), .B2(_0556_ ), .ZN(_0557_ ) );
NAND2_X1 _1238_ ( .A1(_0557_ ), .A2(_0192_ ), .ZN(_0558_ ) );
AOI21_X1 _1239_ ( .A(_0558_ ), .B1(_0035_ ), .B2(_0479_ ), .ZN(_0559_ ) );
NOR3_X1 _1240_ ( .A1(_0133_ ), .A2(_0035_ ), .A3(_0494_ ), .ZN(_0560_ ) );
NAND2_X1 _1241_ ( .A1(_0111_ ), .A2(_0036_ ), .ZN(_0561_ ) );
AOI21_X1 _1242_ ( .A(_0561_ ), .B1(_0383_ ), .B2(_0384_ ), .ZN(_0562_ ) );
OR3_X1 _1243_ ( .A1(_0559_ ), .A2(_0560_ ), .A3(_0562_ ), .ZN(_0655_ ) );
OAI21_X1 _1244_ ( .A(_0236_ ), .B1(_0330_ ), .B2(fanout_net_5 ), .ZN(_0563_ ) );
NAND3_X1 _1245_ ( .A1(_0563_ ), .A2(_0113_ ), .A3(_0219_ ), .ZN(_0564_ ) );
NOR2_X1 _1246_ ( .A1(_0221_ ), .A2(_0621_ ), .ZN(_0565_ ) );
MUX2_X1 _1247_ ( .A(_0565_ ), .B(_0543_ ), .S(fanout_net_3 ), .Z(_0566_ ) );
NOR2_X1 _1248_ ( .A1(_0566_ ), .A2(fanout_net_5 ), .ZN(_0567_ ) );
AOI21_X1 _1249_ ( .A(_0286_ ), .B1(_0523_ ), .B2(_0524_ ), .ZN(_0568_ ) );
OAI21_X1 _1250_ ( .A(_0198_ ), .B1(_0567_ ), .B2(_0568_ ), .ZN(_0569_ ) );
NAND2_X1 _1251_ ( .A1(_0569_ ), .A2(_0192_ ), .ZN(_0570_ ) );
AOI21_X1 _1252_ ( .A(_0198_ ), .B1(_0488_ ), .B2(_0489_ ), .ZN(_0571_ ) );
OAI221_X1 _1253_ ( .A(_0564_ ), .B1(_0398_ ), .B2(_0561_ ), .C1(_0570_ ), .C2(_0571_ ), .ZN(_0656_ ) );
OR3_X1 _1254_ ( .A1(_0254_ ), .A2(_0035_ ), .A3(_0494_ ), .ZN(_0572_ ) );
NOR3_X1 _1255_ ( .A1(_0135_ ), .A2(_0097_ ), .A3(_0119_ ), .ZN(_0573_ ) );
NOR3_X1 _1256_ ( .A1(_0118_ ), .A2(fanout_net_3 ), .A3(_0122_ ), .ZN(_0574_ ) );
NOR2_X1 _1257_ ( .A1(_0573_ ), .A2(_0574_ ), .ZN(_0575_ ) );
MUX2_X1 _1258_ ( .A(_0536_ ), .B(_0575_ ), .S(_0088_ ), .Z(_0576_ ) );
MUX2_X1 _1259_ ( .A(_0576_ ), .B(_0500_ ), .S(_0035_ ), .Z(_0577_ ) );
OAI221_X1 _1260_ ( .A(_0572_ ), .B1(_0411_ ), .B2(_0561_ ), .C1(_0577_ ), .C2(_0277_ ), .ZN(_0657_ ) );
AOI21_X1 _1261_ ( .A(_0042_ ), .B1(_0508_ ), .B2(_0509_ ), .ZN(_0578_ ) );
OAI211_X2 _1262_ ( .A(_0542_ ), .B(fanout_net_5 ), .C1(_0544_ ), .C2(fanout_net_3 ), .ZN(_0579_ ) );
OR3_X1 _1263_ ( .A1(_0232_ ), .A2(fanout_net_3 ), .A3(_0632_ ), .ZN(_0580_ ) );
OAI211_X4 _1264_ ( .A(_0622_ ), .B(fanout_net_3 ), .C1(_0164_ ), .C2(_0017_ ), .ZN(_0581_ ) );
NAND3_X1 _1265_ ( .A1(_0580_ ), .A2(_0625_ ), .A3(_0581_ ), .ZN(_0582_ ) );
AND3_X2 _1266_ ( .A1(_0579_ ), .A2(_0060_ ), .A3(_0582_ ), .ZN(_0583_ ) );
OR3_X2 _1267_ ( .A1(_0578_ ), .A2(_0036_ ), .A3(_0583_ ), .ZN(_0584_ ) );
NAND2_X1 _1268_ ( .A1(_0424_ ), .A2(_0036_ ), .ZN(_0585_ ) );
NAND3_X1 _1269_ ( .A1(_0584_ ), .A2(_0112_ ), .A3(_0585_ ), .ZN(_0586_ ) );
OAI21_X1 _1270_ ( .A(_0586_ ), .B1(_0494_ ), .B2(_0416_ ), .ZN(_0658_ ) );
NAND2_X1 _1271_ ( .A1(_0437_ ), .A2(_0036_ ), .ZN(_0587_ ) );
OR3_X1 _1272_ ( .A1(_0516_ ), .A2(_0042_ ), .A3(_0519_ ), .ZN(_0588_ ) );
OR3_X1 _1273_ ( .A1(_0118_ ), .A2(_0200_ ), .A3(_0122_ ), .ZN(_0589_ ) );
OR2_X4 _1274_ ( .A1(_0121_ ), .A2(_0126_ ), .ZN(_0590_ ) );
OAI211_X2 _1275_ ( .A(_0589_ ), .B(_0286_ ), .C1(fanout_net_3 ), .C2(_0590_ ), .ZN(_0591_ ) );
NAND3_X1 _1276_ ( .A1(_0553_ ), .A2(_0554_ ), .A3(fanout_net_5 ), .ZN(_0592_ ) );
NAND3_X1 _1277_ ( .A1(_0591_ ), .A2(_0153_ ), .A3(_0592_ ), .ZN(_0593_ ) );
NAND3_X1 _1278_ ( .A1(_0588_ ), .A2(_0071_ ), .A3(_0593_ ), .ZN(_0594_ ) );
NAND3_X1 _1279_ ( .A1(_0587_ ), .A2(_0112_ ), .A3(_0594_ ), .ZN(_0595_ ) );
NOR2_X1 _1280_ ( .A1(_0132_ ), .A2(fanout_net_5 ), .ZN(_0596_ ) );
NAND3_X1 _1281_ ( .A1(_0596_ ), .A2(_0113_ ), .A3(_0219_ ), .ZN(_0597_ ) );
NAND2_X1 _1282_ ( .A1(_0595_ ), .A2(_0597_ ), .ZN(_0659_ ) );
NAND3_X1 _1283_ ( .A1(_0219_ ), .A2(_0441_ ), .A3(_0113_ ), .ZN(_0598_ ) );
NOR2_X1 _1284_ ( .A1(_0566_ ), .A2(_0286_ ), .ZN(_0599_ ) );
NOR3_X1 _1285_ ( .A1(_0631_ ), .A2(_0033_ ), .A3(_0627_ ), .ZN(_0600_ ) );
NOR3_X1 _1286_ ( .A1(_0232_ ), .A2(_0168_ ), .A3(_0632_ ), .ZN(_0601_ ) );
NOR3_X1 _1287_ ( .A1(_0600_ ), .A2(_0601_ ), .A3(fanout_net_5 ), .ZN(_0602_ ) );
OAI21_X1 _1288_ ( .A(_0198_ ), .B1(_0599_ ), .B2(_0602_ ), .ZN(_0603_ ) );
NAND2_X1 _1289_ ( .A1(_0603_ ), .A2(_0192_ ), .ZN(_0604_ ) );
AOI21_X1 _1290_ ( .A(_0198_ ), .B1(_0526_ ), .B2(_0527_ ), .ZN(_0605_ ) );
OAI221_X1 _1291_ ( .A(_0598_ ), .B1(_0604_ ), .B2(_0605_ ), .C1(_0451_ ), .C2(_0561_ ), .ZN(_0661_ ) );
NAND4_X1 _1292_ ( .A1(_0455_ ), .A2(_0070_ ), .A3(_0113_ ), .A4(_0071_ ), .ZN(_0606_ ) );
NAND2_X1 _1293_ ( .A1(_0533_ ), .A2(_0537_ ), .ZN(_0607_ ) );
AOI21_X1 _1294_ ( .A(_0131_ ), .B1(_0032_ ), .B2(_0023_ ), .ZN(_0608_ ) );
MUX2_X2 _1295_ ( .A(_0590_ ), .B(_0608_ ), .S(_0097_ ), .Z(_0609_ ) );
MUX2_X2 _1296_ ( .A(_0575_ ), .B(_0609_ ), .S(_0088_ ), .Z(_0610_ ) );
MUX2_X2 _1297_ ( .A(_0607_ ), .B(_0610_ ), .S(_0153_ ), .Z(_0611_ ) );
OAI221_X1 _1298_ ( .A(_0606_ ), .B1(_0465_ ), .B2(_0561_ ), .C1(_0611_ ), .C2(_0277_ ), .ZN(_0662_ ) );
BUF_X1 _1299_ ( .A(\b[2] ), .Z(_0034_ ) );
BUF_X1 _1300_ ( .A(\b[1] ), .Z(_0033_ ) );
BUF_X1 _1301_ ( .A(\a[0] ), .Z(_0000_ ) );
BUF_X1 _1302_ ( .A(\a[1] ), .Z(_0011_ ) );
BUF_X1 _1303_ ( .A(\b[0] ), .Z(_0032_ ) );
BUF_X1 _1304_ ( .A(\a[2] ), .Z(_0022_ ) );
BUF_X1 _1305_ ( .A(\a[3] ), .Z(_0025_ ) );
BUF_X1 _1306_ ( .A(\a[4] ), .Z(_0026_ ) );
BUF_X1 _1307_ ( .A(\a[5] ), .Z(_0027_ ) );
BUF_X1 _1308_ ( .A(\a[6] ), .Z(_0028_ ) );
BUF_X1 _1309_ ( .A(\a[7] ), .Z(_0029_ ) );
BUF_X1 _1310_ ( .A(\a[8] ), .Z(_0030_ ) );
BUF_X1 _1311_ ( .A(\a[9] ), .Z(_0031_ ) );
BUF_X1 _1312_ ( .A(\a[10] ), .Z(_0001_ ) );
BUF_X1 _1313_ ( .A(\a[11] ), .Z(_0002_ ) );
BUF_X1 _1314_ ( .A(\a[12] ), .Z(_0003_ ) );
BUF_X1 _1315_ ( .A(\a[13] ), .Z(_0004_ ) );
BUF_X1 _1316_ ( .A(\a[14] ), .Z(_0005_ ) );
BUF_X1 _1317_ ( .A(\a[15] ), .Z(_0006_ ) );
BUF_X1 _1318_ ( .A(\b[3] ), .Z(_0035_ ) );
BUF_X1 _1319_ ( .A(\a[16] ), .Z(_0007_ ) );
BUF_X1 _1320_ ( .A(\a[17] ), .Z(_0008_ ) );
BUF_X1 _1321_ ( .A(\a[18] ), .Z(_0009_ ) );
BUF_X1 _1322_ ( .A(\a[19] ), .Z(_0010_ ) );
BUF_X1 _1323_ ( .A(\a[20] ), .Z(_0012_ ) );
BUF_X1 _1324_ ( .A(\a[21] ), .Z(_0013_ ) );
BUF_X1 _1325_ ( .A(\a[22] ), .Z(_0014_ ) );
BUF_X1 _1326_ ( .A(\a[23] ), .Z(_0015_ ) );
BUF_X1 _1327_ ( .A(\a[24] ), .Z(_0016_ ) );
BUF_X1 _1328_ ( .A(\a[25] ), .Z(_0017_ ) );
BUF_X1 _1329_ ( .A(\a[26] ), .Z(_0018_ ) );
BUF_X1 _1330_ ( .A(\a[27] ), .Z(_0019_ ) );
BUF_X1 _1331_ ( .A(\a[28] ), .Z(_0020_ ) );
BUF_X1 _1332_ ( .A(\a[29] ), .Z(_0021_ ) );
BUF_X1 _1333_ ( .A(\a[30] ), .Z(_0023_ ) );
BUF_X1 _1334_ ( .A(\a[31] ), .Z(_0024_ ) );
BUF_X1 _1335_ ( .A(\b[4] ), .Z(_0036_ ) );
BUF_X1 _1336_ ( .A(\ctrl[1] ), .Z(_0038_ ) );
BUF_X1 _1337_ ( .A(\ctrl[0] ), .Z(_0037_ ) );
BUF_X1 _1338_ ( .A(\ctrl[3] ), .Z(_0040_ ) );
BUF_X1 _1339_ ( .A(\ctrl[2] ), .Z(_0039_ ) );
BUF_X1 _1340_ ( .A(_0638_ ), .Z(\result[0] ) );
BUF_X1 _1341_ ( .A(_0649_ ), .Z(\result[1] ) );
BUF_X1 _1342_ ( .A(_0660_ ), .Z(\result[2] ) );
BUF_X1 _1343_ ( .A(_0663_ ), .Z(\result[3] ) );
BUF_X1 _1344_ ( .A(_0664_ ), .Z(\result[4] ) );
BUF_X1 _1345_ ( .A(_0665_ ), .Z(\result[5] ) );
BUF_X1 _1346_ ( .A(_0666_ ), .Z(\result[6] ) );
BUF_X1 _1347_ ( .A(_0667_ ), .Z(\result[7] ) );
BUF_X1 _1348_ ( .A(_0668_ ), .Z(\result[8] ) );
BUF_X1 _1349_ ( .A(_0669_ ), .Z(\result[9] ) );
BUF_X1 _1350_ ( .A(_0639_ ), .Z(\result[10] ) );
BUF_X1 _1351_ ( .A(_0640_ ), .Z(\result[11] ) );
BUF_X1 _1352_ ( .A(_0641_ ), .Z(\result[12] ) );
BUF_X1 _1353_ ( .A(_0642_ ), .Z(\result[13] ) );
BUF_X1 _1354_ ( .A(_0643_ ), .Z(\result[14] ) );
BUF_X1 _1355_ ( .A(_0644_ ), .Z(\result[15] ) );
BUF_X1 _1356_ ( .A(_0645_ ), .Z(\result[16] ) );
BUF_X1 _1357_ ( .A(_0646_ ), .Z(\result[17] ) );
BUF_X1 _1358_ ( .A(_0647_ ), .Z(\result[18] ) );
BUF_X1 _1359_ ( .A(_0648_ ), .Z(\result[19] ) );
BUF_X1 _1360_ ( .A(_0650_ ), .Z(\result[20] ) );
BUF_X1 _1361_ ( .A(_0651_ ), .Z(\result[21] ) );
BUF_X1 _1362_ ( .A(_0652_ ), .Z(\result[22] ) );
BUF_X1 _1363_ ( .A(_0653_ ), .Z(\result[23] ) );
BUF_X1 _1364_ ( .A(_0654_ ), .Z(\result[24] ) );
BUF_X1 _1365_ ( .A(_0655_ ), .Z(\result[25] ) );
BUF_X1 _1366_ ( .A(_0656_ ), .Z(\result[26] ) );
BUF_X1 _1367_ ( .A(_0657_ ), .Z(\result[27] ) );
BUF_X1 _1368_ ( .A(_0658_ ), .Z(\result[28] ) );
BUF_X1 _1369_ ( .A(_0659_ ), .Z(\result[29] ) );
BUF_X1 _1370_ ( .A(_0661_ ), .Z(\result[30] ) );
BUF_X1 _1371_ ( .A(_0662_ ), .Z(\result[31] ) );
BUF_X8 fanout_buf_1 ( .A(_0032_ ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(_0033_ ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(_0033_ ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(_0034_ ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(_0034_ ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(_0035_ ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(_0036_ ), .Z(fanout_net_7 ) );

endmodule
