`include "../inc/defines.svh"

module pmu (

);

endmodule